f<int> main() {
    // Plus
    printf("Result: %s\n", String("Hello ") + String("World!"));
    String s1 = String("Hello ") + String("World!");
    printf("Result: %s\n", s1);
    printf("Result: %s\n", s1 + " Hi!");
    printf("Result: %s\n", String("Hi! ") + s1);
    printf("Result: %s\n", s1 + s1);
    printf("Result: %s\n", s1 + " " + s1);
    printf("Result: %s\n", String("Prefix ") + s1 + " Suffix");

    // Mul
    printf("Result: %s\n", 4s * String("Hi"));
    String s2 = String("Hello ") * 5;
    printf("Result: %s\n", s2);
    printf("Result: %s\n", 20 * String('a'));
    String s3 = 2 * String('c') * 7;
    printf("Result: %s\n", s3);

    // Equals raw
    printf("Equal: %d\n", "Hello World!" == "Hello Programmers!");
    printf("Equal: %d\n", "Hello" == "Hell2");
    printf("Equal: %d\n", "Hello" == "Hello");

    // Equals
    printf("Equal: %d\n", String("Hello World!") == String("Hello Programmers!"));
    printf("Equal: %d\n", String("Hello") == String("Hell2"));
    printf("Equal: %d\n", String("Hello") == String("Hello"));

    // Not equals raw
    printf("Non-equal: %d\n", "Hello World!" != "Hello Programmers!");
    printf("Non-equal: %d\n", "Hello" != "Hell2");
    printf("Non-equal: %d\n", "Hello" != "Hello");

    // Not equals
    printf("Non-equal: %d\n", String("Hello World!") != String("Hello Programmers!"));
    printf("Non-equal: %d\n", String("Hello") != String("Hell2"));
    printf("Non-equal: %d\n", String("Hello") != String("Hello"));

    // PlusEquals
    String s4 = String("Hello");
    s4 += 'l';
    printf("Result: %s\n", s4);
    String s5 = String("Hi");
    s5 += " World!";
    printf("Result: %s\n", s5);

    // MulEquals
    String s6 = String("Hi");
    s6 *= 3;
    printf("Result: %s\n", s6);
}