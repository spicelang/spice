type T dyn;

f<int> main() {
    printf("Size: %d", sizeof(T));
}