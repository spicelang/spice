type Alias alias int;
type Alias alias double;

f<int> main() {}