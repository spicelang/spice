import "std/text/print" as print;

type Test struct {
    int field1
    byte field2
}

f<int> Test.getField1() {
    return this.field1;
}

p Test.print(bool b) {
    if b {
        printf("Content: %d, %d", this.field1, this.field2);
    }
}

f<int> main() {
    byte b = 50;
    Test test = new Test { 1, b };
    int field1 = test.getField1();
    printf("Field1: %d", field1);
    print.println("Test");
    //test.print();
}