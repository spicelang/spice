import "std/io/dir" as dir;

f<int> main() {
    printf("Existing before create: %d\n", dir.dirExists("./test"));
    dyn mkReturnCode = dir.mkDir("./test", dir.MODE_ALL_RWX);
    printf("mkDir return code: %d\n", mkReturnCode);
    printf("Existing after create: %d\n", dir.dirExists("./test"));
    dyn rmReturnCode = dir.rmDir("./test");
    printf("rmDir return code: %d\n", rmReturnCode);
    printf("Existing after delete: %d\n", dir.dirExists("./test"));
}