f<double> calledFunction(int mandatoryArg, dyn optionalArg = true) {
    printf("Mandatory: %d", mandatoryArg);
    printf("Optional: %d", optionalArg);
    return 0.1;
}

f<double> calledFunction(string testString) {
    printf("String: %s", testString);
    return 0.3;
}

f<int> main() {
    dyn res = calledFunction(1, false);
    printf("Result: %f", res);
    calledFunction("test");
}