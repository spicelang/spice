f<int> main() {
    short s = 123s;
    dyn** dynPointer = &&s;
}