import "source3" as s3;

public f<int> forwardToOtherModule() {
    result = s3::spawnInteger();
    printf("Spawned integer: %d", result);
}