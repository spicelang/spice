f<int> main() {
    short s = 10;
    s = s + 1;
    long l = 10;
    printf("Short: %d, Long: %d\n", s, l);
}