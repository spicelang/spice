/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = new StringStruct {};
    a.appendChar('A');
}*/

import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = new str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}