/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

f<int> makePi() {
    // Initialize variables
    int q = 1;
    int r = 0;
    int t = 1;
    int k = 1;
    int m = 3;
    int x = 3;
    // Loop
    //int[1000] output = {};
    int outputCounter = 0;
    for int i = 0; i < 1000; i++ {
        if (4 * q + r - t < m * t) {
            //output[outputCounter] = m;
            outputCounter++;
            q = 10 * q;
            r = 10 * (r - m * t);
            t = t;
            k = k;
            m = (10 * (3 * q + r)) / t - 10 * m;
            x = x;
        } else {
            q = q * k;
            r = (2 * q + r) * x;
            t = t * x;
            k = k + 1;
            m = (q * (7 * k + 2) + r * x) / (t * x);
            x = x + 2;
        }
    }
    return 3;
}

f<int> main() {
    makePi();
}