import "std/os/thread";

ext p usleep(int);

p threadRoutine() {
    printf("Test\n");
    printf("Hello from thread: %d\n", getThreadId());
}

f<int> main() {
    Thread t1 = Thread(threadRoutine);
    Thread t2 = Thread(threadRoutine);
    t1.join();
    t2.join();
}