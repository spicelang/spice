public type IStruct interface {

}
