import "std/io/file" as file;

f<int> main() {
    file.FilePtr fp = file.openFile("./test.txt", file.MODE_WRITE);
    fp.writeChar('A');
    fp.close();
}