// Imports
import "std/type/string" as str;

// Constants
const unsigned long INITIAL_ALLOC_COUNT = 5l;
const unsigned int RESIZE_FACTOR = 2;

// Link external functions
ext<byte*> malloc(long);
ext<byte*> realloc(byte*, int);
ext free(byte*);
ext<byte*> memcpy(byte*, byte*, int);

/**
 * String wrapper for enriching raw strings with information and make them mutable
 */
public type String struct {
    char* contents         // Pointer to the first char
    unsigned long capacity // Allocated number of chars
    unsigned long length   // Current number of chars
}

public p String.ctor(const string value = "") {
    this.length = str.getRawLength(value);
    this.capacity = this.length > INITIAL_ALLOC_COUNT ? this.length * RESIZE_FACTOR : INITIAL_ALLOC_COUNT; // +1 because of null terminator

    // Allocate space for the initial number of elements
    unsafe {
        this.contents = (char*) malloc(sizeof(type char) * this.capacity);
    }

    // Save initial value
    unsafe {
        for unsigned long i; i < this.length + 1; i++ { // +1 because of null terminator
            this.contents[i] = value[i];
        }
    }
}

public p String.ctor(const string value1, const string value2) {
    unsigned long value1Length = str.getRawLength(value1);
    unsigned long value2Length = str.getRawLength(value2);
    this.length = value1Length + value2Length;
    this.capacity = this.length > INITIAL_ALLOC_COUNT ? this.length * RESIZE_FACTOR : INITIAL_ALLOC_COUNT; // +1 because of null terminator

    // Allocate space for the initial number of elements
    unsafe {
        this.contents = (char*) malloc(sizeof(type char) * this.capacity);
    }

    // Save initial value
    unsafe {
        for unsigned long i; i < value1Length; i++ {
            this.contents[i] = value1[i];
        }
        for unsigned long i; i < value2Length + 1; i++ { // +1 because of null terminator
            this.contents[value1Length + i] = value2[i];
        }
    }
}

public p String.ctor(const char value) {
    this.length = 1l;
    this.capacity = INITIAL_ALLOC_COUNT;

    // Allocate space for the initial number of elements
    unsafe {
        this.contents = (char*) malloc(sizeof(type char) * this.capacity);
    }

    // Save initial value
    unsafe {
        this.contents[0] = value;
        this.contents[1] = '\0';
    }
}

public p String.dtor() {
    // Free all the memory
    unsafe {
        free((byte*) this.contents);
    }
}

/**
 * Appends the given string wrapper to the current one
 *
 * @param appendix string to be appended
 */
public p String.append(const string appendix) {
    unsigned long appendixLength = str.getRawLength(appendix);
    // Check if we need to re-allocate memory
    while this.capacity <= this.length + appendixLength {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Save data
    unsafe {
        for int i = 0; i < appendixLength + 1; i++ { // +1 because of null terminator
            this.contents[this.length++] = appendix[i];
        }
    }
    this.length--; // Remove null terminator
}

/**
 * Appends the given char to the string and resize it if needed
 *
 * @param c Char to append
 */
public p String.append(const char c) {
    // Check if we need to re-allocate memory
    if this.capacity <= this.length + 1 {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Insert the char at the right position
    unsafe {
        this.contents[this.length++] = c;
        this.contents[this.length] = '\0';
    }
}

/**
 * Implements the multily operator for 'string * int' or 'int * string'
 *
 * @param operand Number of repetitions
 */
public inline p String.opMul(const int operand) {
    this.opMul((long) operand);
}

/**
 * Implements the multily operator for 'string * long' or 'long * string'
 *
 * @param operand Number of repetitions
 */
public p String.opMul(const long operand) {
    // Cancel if operand is less than 2
    if operand < 2l { return; }

    unsigned long newLength = operand * this.length;
    // Check if we need to re-allocate memory
    while this.capacity <= newLength {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Save the value
    unsafe {
        for unsigned long i = 0l; i < newLength; i++ {
            this.contents[i] = this.contents[i % this.length];
        }
        this.contents[newLength] = '\0';
    }
    this.length = newLength;
}

/**
 * Implements the multily operator for 'string * short' or 'short * string'
 *
 * @param operand Number of repetitions
 */
public inline p String.opMul(const short operand) {
    this.opMul((long) operand);
}

/**
 * Implements the equals operator for 'string == string'
 *
 * @param operand String to comare the current string to
 *
 * @return Equal or not
 */
public f<bool> String.opEquals(const string operand) {
    // Compare sizes
    if str.getRawLength(operand) != this.length {
        return false;
    }

    // Compare contents
    unsafe {
        for int i = 0; i < this.length; i++ {
            if this.contents[i] != operand[i] {
                return false;
            }
        }
    }

    return true;
}

/**
 * Implements the equals operator for 'string != string'
 *
 * @param operand String to comare the current string to
 *
 * @return Equal or not
 */
public inline f<bool> String.opNotEquals(const string operand) {
    return !this.opEquals(operand);
}

/**
 * Get the raw and immutable string from this container instance
 *
 * @return Raw immutable string
 */
public inline f<string> String.getRaw() {
    return (string) this.contents;
}

/**
 * Retrieve the current length of the string
 *
 * @return Current length of the string
 */
public inline f<long> String.getLength() {
    return this.length;
}

/**
 * Check if the string is empty
 */
public inline f<bool> String.isEmpty() {
    return this.length == 0;
}

/**
 * Retrieve the current capacity of the string
 *
 * @return Current capacity of the string
 */
 public inline f<long> String.getCapacity() {
     return this.capacity - 1; // -1 because of null terminator
 }

/**
 * Checks if the string exhausts its capacity
 *
 * @return Full or not full
 */
public inline f<bool> String.isFull() {
    return this.length == this.capacity;
}

/**
 * Replaces the current contents of the string with an empty string
 */
public p String.clear() {
    this.length = 0l;
    unsafe {
        this.contents[0] = '\0';
    }
}

/**
 * Reserves `charCount` items
 *
 * @param charCount Number of chars to reserve for the string
 */
public p String.reserve(unsigned long charCount) {
    if charCount > this.capacity {
        this.resize(charCount);
    }
}

/**
 * Re-allocates heap space for the string contents
 *
 * @param newLength new length of the string after resizing
 */
p String.resize(unsigned long newLength) {
    // Allocate the new memory
    unsafe {
        byte* oldAddress = (byte*) this.contents;
        int newSize = (int) (sizeof(type char) * newLength);
        char* newMemory = (char*) realloc(oldAddress, newSize);
        this.contents = newMemory;
    }
    // Set new capacity
    this.capacity = newLength;
}