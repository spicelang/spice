f<int> add(int a, int b) {
    return a + b;
}

#[test]
f<bool> testAdd() {
    assert add(1, 2) == 4; // Failing assertion means the test failed
    return true;
}
