// Imports
import "std/type/type-conversion";

public type CodeLoc struct {
    public unsigned long line
    public unsigned long col
    public string sourceFilePath
}

public p CodeLoc.ctor(unsigned long line, unsigned long col, string sourceFilePath = "") {
    this.line = line;
    this.col = col;
    this.sourceFilePath = sourceFilePath;
}

/**
 * Returns the code location as a string for using it as a map key or similar
 *
 * @return Code location string
 */
public f<String> CodeLoc.toString() {
    return "L" + toString(this.line) + "C" + toString(this.col);
}

/**
 * Returns the code location in a pretty form
 *
 * @return Pretty code location
 */
public f<String> CodeLoc.toPrettyString() {
    if len(this.sourceFilePath) == 0 {
        return toString(this.line) + ":" + toString(this.col);
    }
    return this.sourceFilePath + ":" + toString(this.line) + ":" + toString(this.col);
}

/**
 * Returns the line number in a pretty form
 *
 * @return Pretty line number
 */
public f<String> CodeLoc.toPrettyLine() {
    return "L" + toString(this.line);
}

/**
 * Returns the line and column number in a pretty form
 */
public f<String> CodeLoc.toPrettyLineAndColumn() {
    return this.toString();
}

public f<bool> operator==(const CodeLoc &lhs, const CodeLoc &rhs) {
    return lhs.sourceFilePath == rhs.sourceFilePath && lhs.line == rhs.line && lhs.col == rhs.col;
}