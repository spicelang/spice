import "std/data/red-black-tree";
import "std/iterator/iterable";
import "std/iterator/iterator";
import "std/data/pair";

// Add generic type definitions
type K dyn;
type V dyn;

/**
 * A map in Spice is a commonly used data structure, which can be used to represent a list of key value pairs.
 *
 * Time complexity:
 * Insert: O(log n)
 * Delete: O(log n)
 * Lookup: O(log n)
 */
public type Map<K, V> struct : IIterable<Pair<K, V>> {
    RedBlackTree<K, V> tree
}

/**
 * Inserts a key value pair into the map.
 *
 * @param key The key to insert.
 * @param value The value to insert.
 */
public p Map.insert(const K& key, const V& value) {
    this.tree.insert(key, value);
}

/**
 * Removes a key value pair from the map.
 *
 * @param key The key to remove.
 */
public p Map.remove(const K& key) {
    this.tree.remove(key);
}

/**
 * Retrieve the value associated with the given key.
 * Note: If the key is not found in the map, this function will panic. To avoid this, use getSafe instead.
 *
 * @param key The key to get.
 * @return The value associated with the key.
 */
public f<V&> Map.get(const K& key) {
    return this.tree.find(key);
}

/**
 * Retrieve the value associated with the given key.
 * Note: If the key is not found in the map, this function will panic. To avoid this, use getSafe instead.
 *
 * @param key The key to get.
 * @return The value associated with the key.
 */
public f<V&> operator[]<K, V>(Map<K, V>& map, const K& key) {
    return map.get(key);
}

/**
 * Retrieve the value associated with the given key as Result<V>.
 * If the key is not found, the result contains an error.
 *
 * @param key The key to look up
 * @return Result<V>, containing the value associated with the key or an error if the key is not found
 */
public f<Result<V>> Map.getSafe(const K& key) {
    return this.tree.findSafe(key);
}

/**
 * Checks if the map contains a key.
 *
 * @param key The key to check.
 * @return True if the map contains the key, false otherwise.
 */
public f<bool> Map.contains(const K& key) {
    return this.tree.contains(key);
}

/**
 * Gets the number of elements in the map.
 *
 * @return The number of elements in the map.
 */
public f<unsigned long> Map.getSize() {
    return this.tree.getSize();
}

/**
 * Checks if the map is empty.
 *
 * @return True if the map is empty, false otherwise.
 */
public f<bool> Map.isEmpty() {
    return this.tree.getSize() == 0l;
}

/**
 * Removes all elements from the map.
 */
public p Map.clear() {
    this.tree.clear();
}

/**
 * Iterator to iterate over a map data structure
 */
public type MapIterator<K, V> struct : IIterator<Pair<const K&, V&>> {
    RedBlackTreeIterator<K, V> rbtIterator
}

public p MapIterator.ctor<K, V>(Map<K, V>& map) {
    this.rbtIterator = map.tree.getIterator();
}

/**
 * Returns the current key-value pair of the map
 *
 * @return Current key/value pair
 */
public inline f<Pair<const K&, V&>&> MapIterator.get() {
    return this.rbtIterator.get();
}

/**
 * Returns the current index and the current item of the map
 *
 * @return Pair of current index and current key/value pair
 */
public inline f<Pair<unsigned long, Pair<const K&, V&>&>> MapIterator.getIdx() {
    return this.rbtIterator.getIdx();
}

/**
 * Check if the iterator is valid
 *
 * @return true or false
 */
public inline f<bool> MapIterator.isValid() {
    return this.rbtIterator.isValid();
}

/**
 * Moves the cursor to the next key/value pair
 */
public inline p MapIterator.next() {
    this.rbtIterator.next();
}

/**
 * Advances the cursor by one
 *
 * @param it MapIterator
 */
public inline p operator++<K, V>(MapIterator<K, V>& it) {
    this.htIterator.next();
}

/**
 * Retrieve a forward iterator for the map
 */
public f<MapIterator<K, V>> Map.getIterator() {
    return MapIterator<K, V>(*this);
}
