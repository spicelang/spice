// Imports

public type EntryNode struct {

}