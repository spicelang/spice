// Link external functions
ext f<heap byte*> malloc(long);
ext p free(heap byte*);

// Add generic type definitions
type T dyn;

// Enums
type NodeColor enum { RED, BLACK }

/**
 * Node of a Red-Black Tree
 */
type Node<T> struct {
    T data
    heap Node<T>* childLeft
    heap Node<T>* childRight
    NodeColor color
}

f<Node<T>*> createNode<T>(T data) {
    heap Node<T>* newNode = (heap Node<T>*) malloc(sizeof(type Node<T>) / 8);
    newNode.data = data;
    newNode.childLeft = nil<heap Node<T>*>;
    newNode.childRight = nil<heap Node<T>*>;
    newNode.color = NodeColor::RED;
    return newNode;
}

inline f<bool> Node.isRoot() {
    return this.parent == nil<heap Node<T>*>;
}

/**
 * A Red-Black Tree is a self-balancing search tree, which is used e.g. in the implementation of maps.
 *
 * Insertion time: O(log n)
 * Lookup time: O(log n)
 * Deletion time: O(log n)
 */
public type RedBlackTree<T> struct {
    heap Node<T>* rootNode
}

public p RedBlackTree.ctor() {
    this.rootNode = nil<heap Node<T>*>;
}

public p RedBlackTree.insert(T newItem) {
    this.insertAdd(newItem);
    this.insertRebalance(newItem);
}

p RedBlackTree.insertAdd(T newItem) {

}

p RedBlackTree.insertRebalance(T newItem) {

}