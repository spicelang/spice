type Result struct {}

f<int> main() {
    Result res;
}