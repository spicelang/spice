import "std/iterator/number-iterator";

f<int> main() {
    dyn shortIterator = range(3s, 8s);
    foreach short s : shortIterator {
        printf("Short %d\n", s);
        if ((s & 1s) == 1) {
            foreach dyn l : range(1l, 2l) {
                printf("Long %d\n", l);
                break 2;
            }
        }
    }
    printf("End.");
}