import "test2" as s1;

f<int> main() {
    dyn v = s1::Vector<int>{};
    v.setData(12);
    printf("Data: %d\n", v.data);
    v.setData(1.5);
    printf("Data: %d\n", v.data);
}

/*import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

public type TestNode struct {
    int data = 123
}

public p TestNode.dtor() {}

f<int> main() {
    DefaultMemoryManager mm;
    BlockAllocator<TestNode> ba = BlockAllocator<TestNode>(mm);
}*/