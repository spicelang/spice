import "std/type/result";

f<int> main() {
    Result<int> r = ok(1);
    printf("%d", r.unwrap());
}

/*type A struct {
    int f1
}

type B struct {
    int f3
}

type C struct {
    compose A _1
    compose B _2
    int f2
}

f<int> main() {
    C c;
    c.f1 = 1;
    c.f2 = 2;
    c.f3 = 3;
    printf("%d, %d, %d\n", c.f1, c.f2, c.f3);
}*/