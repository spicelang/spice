type T dyn;

f<int> print<T>(T g) {
    printf("%d", g);
    return 0;
}

f<int> main() {
    print(1);
    print("string");
}