public type IScope interface {

}
