/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec.Vector<pair.Pair<int, string>> pairVector = vec.Vector<pair.Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair.Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

type TestStruct struct {
    bool test
}

p TestStruct.dtor(int test) {
    printf("Dtor called");
}

f<int> main() {
    TestStruct t = TestStruct();
    printf("Test: %d\n", 0o0000777);
}