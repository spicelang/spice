f<int> malloc(int size) {
    // ToDo: Implement @marcauberer
    return 0;
}