f<int> main() {
    const int constVar = 101;
    constVar++;
}