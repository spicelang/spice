f<int> main() {
    printf("Output: %s", test);
    return 0;
}