f<int> main() {
    int arraySize = 4;
    int[arraySize] intArray;
    intArray[1] = 12;
    intArray[2] = 7;
    //printf("Size: %d\n", len(intArray));
}