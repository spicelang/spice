f<int> main() {
    for dyn i = 0; i < 10; i+=2 {
        printf("Step %d\n", i);
    }
}