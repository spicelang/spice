f<int> main() {
    int test = 12;
    int* testPtr = &test;
    printf("Pointer: %p, value: %d", testPtr, test);
}