type T1 dyn;
type T2 dyn;

type Test struct {}

inline f<bool> isSame<T1, T2>() {
    if typeid<T1>() == typeid<T2>() {
        return true;
    } else {
        return false;
    }
}

f<int> main() {
    printf("%d\n", isSame<Test, Test>());
    printf("%d\n", isSame<Test, int>());
    printf("%d\n", isSame<double*, Test>());
}