p foo() {
    panic(Error("This is an error"));
}

f<int> main() {
    foo();
}