/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec::Vector<pair::Pair<int, string>> pairVector = vec.Vector<pair::Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair::Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

import "std/runtime/string_rt" as _rt_str;

f<int> main() {
    // Plus
    printf("Result: %s\n", "Hello " + "World!");
    string s1 = "Hello " + "World!";
    printf("Result: %s\n", s1);
    // Mul
    printf("Result: %s\n", 4s * "Hi");
    string s2 = "Hello " * 5;
    printf("Result: %s\n", s2);
    // Equals
    printf("Equal: %d\n", "Hello World!" == "Hello Programmers!");
    printf("Equal: %d\n", "Hello" == "Hell2");
    printf("Equal: %d\n", "Hello" == "Hello");
    // Not equals
    printf("Non-equal: %d\n", "Hello World!" != "Hello Programmers!");
    printf("Non-equal: %d\n", "Hello" != "Hell2");
    printf("Non-equal: %d\n", "Hello" != "Hello");
    // PlusEquals
    string s3 = "Hello";
    s3 += 'l';
    printf("Result: %s\n", s3);
    string s4 = "Hi";
    s4 += " World!";
    printf("Result: %s\n", s4);
}