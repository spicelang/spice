import "std/type/bool";

f<int> main() {
    printf("Result: %d\n", toInt(true));
}