f<int> main() {
    switch 1 {
        case 1.0: { return 1; }
        default: { return 0; }
    }
}
