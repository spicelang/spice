f<int> main() {

}