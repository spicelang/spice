f<int> main() {
    const int test = 12;
    int& ref = test;
    ref++;
}