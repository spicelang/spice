f<int> main() {
    char c = '\x';
}