type String struct {
    int[] value
    int len // Length of the string
    int cap // Capacity of the string. Is always the next higher power of two than len
}

f<String> create(string input) {
    result.value = input;
    result.len = sizeof(input) * 8;
}

p clear(String* strRef) {
    *strRef.value = "";
    *strRef.len = 0;
}

f<int> len(String* strRef) {
    
}

f<String> concat(String a, String b) {
    // Return b if a is empty
    int aLen = len(a);
    if aLen == 0 { return b; }
    // Return a if b is empty
    int bLen = len(b);
    if bLen == 0 { return a; }
    
    // Create a new string on the heap
    // ToDo @marcauberer

    return "";
}