import "std/type/result";
import "std/type/error";

type FilePtr alias byte*;
public type File struct {
    FilePtr* filePtr
}

// Link external functions
ext f<FilePtr*> fopen(string, string);

public f<Result<File>> openFile(string path, string mode) {
    FilePtr* fp = fopen(path, mode);
    File file = File{fp};
    return fp != nil<FilePtr*> ? ok(file) : err(file, Error("Failed to open file"));
}