type T dyn;
type U int|double;

type Node<T, U> struct {
    T* _data1
    U _data2
}

f<int> main() {
    dyn _node = Node<Node<Node<Node<Node<string, double>, int>, double>, int>, double>{};
}

/*import "std/data/stack";

f<int> main() {
    Stack<int> s1 = Stack<int>{};
    s1.ctor();
    s1.push(123);
    s1.push(456);
    s1.push(789);
    printf("Stack size: %d\n", s1.getSize());
    printf("Stack capacity: %d\n", s1.getCapacity());
    printf("Stack item 3: %d\n", s1.pop());
    printf("Stack item 2: %d\n", s1.pop());
    printf("Stack item 1: %d\n", s1.pop());
}*/

/*type TestStruct struct {
    int a = 123
    short b = 1s
}

f<int> main() {
    TestStruct ts;
    printf("%d %d\n", ts.a, ts.b);
}*/