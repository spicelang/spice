f<bool> equal(int a, int b) {
    return a == b;
}

f<int> main() {
    if equal(1, 2) {
        printf("true");
        return 0;
    }
    printf("false");
}