f<int> fib(int n) {
    if n <= 2 { return 1; }
    return fib(n - 1) + fib(n - 2);
}

f<int> main() {
    int base = 46
    printf("Fibonacci of %d: %d", base, fib(base));
}