#![core.linker.flag = "-pthread"]

ext f<int> pthread_create(long*, byte*, p(), byte*);
ext f<int> pthread_join(long, byte**);

f<int> main() {
    long tid1;
    long tid2;
    int i = 123;
    pthread_create(&tid1, nil<byte*>, p() {
        i++;
        printf("Hello from thread 1\n");
    }, nil<byte*>);
    pthread_create(&tid2, nil<byte*>, p() {
        i++;
        printf("Hello from thread 2\n");
    }, nil<byte*>);
    pthread_join(tid1, nil<byte**>);
    pthread_join(tid2, nil<byte**>);
    printf("%d\n", i);
}

/*f<int> main() {
    int i = 123; // Captured by ref
    int j = 321; // Captured by val
    dyn lambda = p() {
        printf("Hello from inside: %d\n", i);
        i++;
        i += j;
        printf("Hello from inside: %d\n", i);
    };
    lambda();
    printf("Hello from outside: %d\n", i);
}*/

/*type Visitable interface {
    p print();
}

type Test1 struct : Visitable {
    int f1
}

p Test1.print() {
    printf("Foo: %d", this.f1);
}

f<int> main() {
    Test1 t1 = Test1{123};
    Visitable* v = &t1;
    v.print();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";

f<int> main() {
    Lexer lexer = Lexer("./file.spice");
    Parser parser = Parser(lexer);
    parser.parse();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "std/time/timer";

f<int> main() {
    Timer timer = Timer();
    timer.start();
    Lexer lexer = Lexer("./file.spice");
    unsigned long i = 1l;
    while (!lexer.isEOF()) {
        Token token = lexer.getToken();
        //printf("Token %d: ", i);
        //token.print();
        lexer.advance();
        i++;
    }
    timer.stop();
    printf("Tokens: %d, Time: %d\n", i, timer.getDurationInMillis());
}*/