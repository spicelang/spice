// TEST: --output-container=obj

f<int> add(int a, int b) {
    return a + b;
}