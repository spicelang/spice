f<int> main() {
    if false {
        printf("If content!");
    }
    while true {
        printf("While content!");
    }
    /*int i = 0;
    while i < 5 {
        i++;
    }*/
    /*for int i = 0; i < 3; i++ {
        printf("For content!");
    }*/
    printf("Hello World!");
    printf("Dies ist ein Test: %d, %d", 1, 5);
    return 0;
}