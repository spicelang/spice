type T dyn;
type T int|double;

f<int> main() {}