type i32 alias int;

f<int> main() {
    i32 test = 12;
    printf("Hello World: %d\n", test);
}

/*f<int> main() {
    String s = String("Hello ");
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.append("World!");
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.append('?');
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.append('!');
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    printf("Equals: %d\n", s.isEqual(String("Hello World!?!")));
    printf("Equals: %d\n", s.isEqual(String("Hello World!!")));
    s.clear();
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.reserve(100l);
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s = String("");
    printf("Empty: %d\n", s.isEmpty());
    s.append('a');
    printf("Empty: %d", s.isEmpty());
}*/

/*f<int> main() {
    String strA = String("Hello ");
    String strB = String("World!");
    printf("A: %s\n", strA);
    printf("B: %s\n", strB);
    printf("C: %s\n", String("Hello ") + String("World!"));
    String d = String("Hello ") + String("World!");
    printf("D: %s\n", d);
}*/