import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

type ASTNode struct {
    int value
}

public p ASTNode.dtor() {
    printf("Dtor called!");
}

f<int> main() {
    DefaultMemoryManager defaultMemoryManager;
    IMemoryManager* memoryManager = &defaultMemoryManager;
    BlockAllocator<ASTNode> allocator = BlockAllocator<ASTNode>(memoryManager, 10l);
}