f<int> main() {
    int test = 123;
    int& testRef = test;
    printf("%p\n", &test);
    printf("%p\n", &testRef);
    assert &test == &testRef;
}