// Imports
import "std/text/print";
import "std/os/cmd";
import "std/io/cli-parser";
import "std/io/cli-subcommand";
import "std/io/cli-option";

/**
 * Representation of the various cli options
 */
public type CliOptions struct {
    public String mainSourceFile // e.g. main.spice
    public String targetTriple   // In format: <arch><sub>-<vendor>-<sys>-<abi>
    public String targetArch
    public String targetVendor
    public String targetOs
    public bool execute = false
    public bool isNativeTarget = true
    public String cacheDir
    public String outputDir      // Where the object files go. Should always be a temp directory
    public String outputPath     // Where the output binary goes.
    public unsigned short compileJobCount = 0s // O for auto
    public bool ignoreCache = false
    public bool printDebugOutput = false
    public bool dumpCST = false
    public bool dumpAST = false
    public bool dumpIR = false
    public bool dumpAssembly = false
    public bool dumpSymbolTable = false
    public bool enableAstOpt = false
    public short optLevel = 2s // -O0 = 0, -O1 = 1, -O2 = 2, -O3 = 3, -Os = 4, -Oz = 5
    public bool generateDebugInfo = false
    public bool disableVerifier = false
    public bool testMode = false
}

/**
 * Helper class to setup the cli interface and command line parser
 */
public type CliInterface struct {
    CliParser cliParser
    public CliOptions cliOptions
    public bool shouldCompile = false
    public bool shouldInstall = false
    public bool shouldExecute = false
}

public p CliInterface.createInterface() {
    this.cliParser = CliParser("Spice", "Spice programming language");
    this.cliParser.setFooter("(c) Marc Auberer 2021-2023");

    // Add version flag
    this.cliParser.setVersion("Spice version 0.14.3\nbuilt by: GitHub Actions\n\n(c) Marc Auberer 2021-2023");

    // Create sub-commands
    this.addBuildSubcommand();
    this.addRunSubcommand();
    this.addInstallSubcommand();
    this.addUninstallSubcommand();

    // ToDo: extend
}

/**
 * Initialize the cli options based on the input of the user
 */
public p CliInterface.enrich() {
    // Propagate target information
    if this.cliOptions.targetTriple.isEmpty() && this.cliOptions.targetArch.isEmpty() {
        // ToDo: Extend
    }

    // Dump AST, IR and symbol table if all debug output is enabled
    if this.cliOptions.printDebugOutput {
        this.cliOptions.dumpAST = true;
        this.cliOptions.dumpIR = true;
        this.cliOptions.dumpSymbolTable = true;
    }
}

/**
 * Add build subcommand to cli interface
 */
p CliInterface.addBuildSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.createSubcommand("build", "Builds your Spice program and emits an executable");
    subCmd.addAlias("b");

    addCompileSubcommandOptions(subCmd);

    // --target-triple
    CliOption<string>& targetOption = subCmd.addOption("--target", this.cliOptions.targetTriple, "Target triple for the emitted executable (for cross-compiling)");
    targetOption.addAlias("--target-triple");
    targetOption.addAlias("-t");
    // --target-arch
    CliOption<string>& targetArchOption = subCmd.addOption("--target-arch", this.cliOptions.targetArch, "Target arch for emitted executable (for cross-compiling)");
    // --target-vendor
    CliOption<string>& targetVendorOption = subCmd.addOption("--target-vendor", this.cliOptions.targetVendor, "Target vendor for emitted executable (for cross-compiling)");
    // --target-os
    CliOption<string>& targetOsOption = subCmd.addOption("--target-os", this.cliOptions.targetOs, "Target OS for emitted executable (for cross-compiling)");

    // --output
    CliOption<string>& outputOption = subCmd.addOption("--output", this.cliOptions.outputPath, "Set the output file path");
    outputOption.addAlias("-o");
    // --debug-info
    CliOption<bool>& debugInfoOption = subCmd.addOption("--debug-info", this.cliOptions.generateDebugInfo, "Generate debug info");
    debugInfoOption.addAlias("-g");
    // --disable-verifier
    CliOption<bool>& disableVerifierOption = subCmd.addOption("--disable-verifier", this.cliOptions.disableVerifier, "Disable LLVM module and function verification");
}

/**
 * Add run subcommand to cli interface
 */
p CliInterface.addRunSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.createSubcommand("run", "Builds your Spice program and runs it immediately");
    subCmd.addAlias("r");

    addCompileSubcommandOptions(subCmd);

    // --output
    CliOption<string>& outputOption = subCmd.addOption("--output", this.cliOptions.outputPath, "Set the output file path");
    outputOption.addAlias("-o");
    // --debug-info
    CliOption<bool>& debugInfoOption = subCmd.addOption("--debug-info", this.cliOptions.generateDebugInfo, "Generate debug info");
    debugInfoOption.addAlias("-g");
    // --disable-verifier
    CliOption<bool>& disableVerifierOption = subCmd.addOption("--disable-verifier", this.cliOptions.disableVerifier, "Disable LLVM module and function verification");
}

/**
 * Add install subcommand to cli interface
 */
p CliInterface.addInstallSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.createSubcommand("install", "Builds your Spice program and installs it to a directory in the PATH variable");
    subCmd.addAlias("i");

    addCompileSubcommandOptions(subCmd);
}

/**
 * Add uninstall subcommand to cli interface
 */
p CliInterface.addUninstallSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.createSubcommand("uninstall", "Builds your Spice program and runs it immediately");
    subCmd.addAlias("u");

    addCompileSubcommandOptions(subCmd);
}

p CliInterface.addCompileSubcommandOptions(CliSubcommand& subCmd) {
    // --debug-output
    CliOption<bool>& debugOutputFlag = subCmd.addFlag("--debug-output", this.cliOptions.printDebugOutput, "Enable debug output");
    debugOutputFlag.addAlias("-d");
    // --dump-cst
    CliOption<bool>& dumpCstFlag = subCmd.addFlag("--dump-cst", this.cliOptions.dumpCST, "Dump CSTs as serialized string and SVG image");
    dumpCstFlag.addAlias("-cst");
    // --dump-ast
    CliOption<bool>& dumpAstFlag = subCmd.addFlag("--dump-ast", this.cliOptions.dumpAST, "Dump ASTs as serialized string and SVG image");
    dumpAstFlag.addAlias("-ast");
    // --dump-symtab
    CliOption<bool>& dumpSymtabFlag = subCmd.addFlag("--dump-symtab", this.cliOptions.dumpSymbolTable, "Dump serialized symbol tables");
    dumpSymtabFlag.addAlias("-symtab");
    // --dump-ir
    CliOption<bool>& dumpIrFlag = subCmd.addFlag("--dump-ir", this.cliOptions.dumpIR, "Dump LLVM-IR");
    dumpIrFlag.addAlias("-ir");
    // --dump-assembly
    CliOption<bool>& dumpAsmFlag = subCmd.addFlag("--dump-assembly", this.cliOptions.dumpAssembly, "Dump assembly code");
    dumpAsmFlag.addAlias("-asm");
    dumpAsmFlag.addAlias("-s");

    // --jobs
    CliOption<bool>& jobsFlag = subCmd.addFlag("--jobs", this.cliOptions.compileJobCount, "Compile jobs (threads), used for compilation");
    jobsFlag.addAlias("-j");
    // --ignore-cache
    subCmd.addFlag("--ignore-cache", this.cliOptions.ignoreCache, "Force re-compilation of all source files");
    // --enable-ast-opt
    subCmd.addFlag("--enable-ast-opt", this.cliOptions.enableAstOpt, "Enable first order optimizations on the AST");

    // Opt levels
    //subCmd.addFlag("-O0", [&]() { this.cliOptions.optLevel = 0; }, "Disable optimization for the output executable.");
    //subCmd.addFlag("-O1", [&]() { this.cliOptions.optLevel = 1; }, "Optimization level 1. Only basic optimization is executed.");
    //subCmd.addFlag("-O2", [&]() { this.cliOptions.optLevel = 2; }, "Optimization level 2. More advanced optimization is applied.");
    //subCmd.addFlag("-O3", [&]() { this.cliOptions.optLevel = 3; }, "Optimization level 3. Aggressive optimization for best performance.");
    //subCmd.addFlag("-Os", [&]() { this.cliOptions.optLevel = 4; }, "Optimization level s. Size optimization for output executable.");
    //subCmd.addFlag("-Oz", [&]() { this.cliOptions.optLevel = 5; }, "Optimization level z. Aggressive optimization for best size.");

    CliOption<string>& fileOption = subCmd.addOption("<main-source-file>", this.cliOptions.mainSourceFile, "MainSourceFile");
    fileOption.setRequired();
    fileOption.check(CliOption::EXISTING_FILE);
}

/**
 * Start the parsing process
 *
 * @param argc Argument count
 * @param argv Argument vector
 * @return Return code
 */
public f<int> CliInterface.parse(int argc, string[] argv) {
    return this.cliParser.parse(argc, argv);
}