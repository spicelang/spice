f<int> main() {
    double calcResult = "No bool" ? 5.6 : 1.0;
}