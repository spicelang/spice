import "std/math/fct" as fct;

f<int> main() {
    printf("Abs (int): %d\n", fct.abs(123));
    printf("Abs (int): %d\n", fct.abs(-137));
    printf("Abs (short): %d\n", fct.abs(56s));
    printf("Abs (short): %d\n", fct.abs(-3s));
    printf("Abs (long): %d\n", fct.abs(1234567890l));
    printf("Abs (long): %d\n", fct.abs(-987654321l));
    printf("Abs (double): %f\n", fct.abs(56.123));
    printf("Abs (double): %f\n", fct.abs(-348.12));

    printf("Cos (int): %d\n", fct.cos(23));
    printf("Cos (short): %d\n", fct.cos(68s));
    printf("Cos (long): %d\n", fct.cos(359l));
}

/*type Visitor struct {

}

type SymbolTable struct {

}

type VisitableNode interface {
    f<bool> accept(Visitor*)
}

type AstNode struct : VisitableNode {

}

f<bool> AstNode.accept(Visitor* v) {
    return true;
}

type AstEntryNode struct : VisitableNode {
    AstNode astNode
    SymbolTable* fctScope
    bool hasArgs
}

f<bool> AstEntryNode.accept(Visitor* v) {
    return true;
}

f<int> main() {
    dyn entryNode = AstEntryNode{};
    printf("%d", entryNode.hasArgs);
}*/

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

/*public f<bool> src(bool x, bool y) {
    return ((x ? 1 : 4) & (y ? 1 : 4)) == 0;
}

public f<int> tgt(int x, int y) {
    return x ^ y;
}

f<int> main() {
    printf("Result: %d, %d", src(false, true), tgt(0, 1));
}*/