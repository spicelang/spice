ext<int> mkdir(char*, byte);

f<int> createDir(char* path, byte mode) {
    return mkdir(path, mode);
}