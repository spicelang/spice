type T double|string;
type TestAlias alias UnknownStruct<T>;

f<int> main() {}