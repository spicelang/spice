import "std/time/delay" as delay;
import "std/os/cpu" as cpu;

type Mutex struct {
	bool occupied
}

/**
 * Acquire the mutex
 */
p Mutex.acquire() {
	while this.occupied {
		cpu.yield();
	}
	this.occupied = true;
}

/**
 * Release the mutex
 */
p Mutex.release() {
	this.occupied = false;
}