type NestedStruct struct {
    double* test
}

type TestStruct struct {
    double f1
    NestedStruct* f2
}

f<int> main() {
    dyn test = 1.2;
    dyn ns = NestedStruct{ &test };
    dyn s = TestStruct{ 5.4, &ns };
    printf("Double: %f\n", *s.f2.test);
}