public f<int> dummy() {
    return 1;
}