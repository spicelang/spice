import "std/data/map";

f<int> main() {
    Map<int, string> map;
}

/*import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

f<int> main() {
    DefaultMemoryManager defaultMemoryManager;
    IMemoryManager* memoryManager = &defaultMemoryManager;
    BlockAllocator<int> allocator = BlockAllocator<int>(memoryManager, 10);
}*/