f<int> main() {
    int calcResult1 = true * "test";
    double calcResult2 = false / 3.90;
    string calcResult3 = true / 4;
    bool calcResult4 = true * false;
}