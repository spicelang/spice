type Person struct {
	string firstName
	string lastName
	int age
}

f<int> main() {
	Person john = Person { "John", "Doe", 46 };
	john.age = 47;
	printf("John's age: %d", john.age);
}