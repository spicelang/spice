/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

f<int> faculty(int input) {
    if input < 2 {
        return 1;
    }
    result = input * faculty(input - 1);
}

f<int> main() {
    dyn input = 10;
    int faculty = faculty(input);
    printf("Faculty of %d is: %d", input, faculty);
}