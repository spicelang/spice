f<int> main() {
    int val = 1;
    val += ((1++)--) * 2 << 2;
    assert val == 9;

    printf("All assertions passed!");
}