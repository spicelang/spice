import "std/math/fct" as fct;

f<int> main() {
    printf("Abs (int): %d\n", fct::abs(123));
    printf("Abs (int): %d\n", fct::abs(-137));
    printf("Abs (short): %d\n", fct::abs(56s));
    printf("Abs (short): %d\n", fct::abs(-3s));
    printf("Abs (long): %lld\n", fct::abs(1234567890l));
    printf("Abs (long): %lld\n", fct::abs(-987654321l));
    printf("Abs (double): %f\n", fct::abs(56.123));
    printf("Abs (double): %f\n", fct::abs(-348.12));

    printf("Max (int, int): %d\n", max(1, 2));
    printf("Max (int, int): %d\n", max(-1, -2));
    printf("Max (short, short): %d\n", max(165s, 263s));
    printf("Max (short, short): %d\n", max(-165s, -263s));
    printf("Max (long, long): %lld\n", max(3495872345l, 239458723l));
    printf("Max (long, long): %lld\n", max(-3495872345l, -239458723l));
    printf("Max (double, double): %f\n", max(34.234971, 34.23497));
    printf("Max (double, double): %f\n", max(-34.234971, -34.23497));

    printf("Min (int, int): %d\n", min(1, 2));
    printf("Min (int, int): %d\n", min(-1, -2));
    printf("Min (short, short): %d\n", min(165s, 263s));
    printf("Min (short, short): %d\n", min(-165s, -263s));
    printf("Min (long, long): %lld\n", min(3495872345l, 239458723l));
    printf("Min (long, long): %lld\n", min(-3495872345l, -239458723l));
    printf("Min (double, double): %f\n", min(34.234971, 34.23497));
    printf("Min (double, double): %f\n", min(-34.234971, -34.23497));

    printf("Trunc (double): %d\n", trunc(1.499));
    printf("Trunc (double): %d\n", trunc(1.500));
    printf("Trunc (double): %d\n", trunc(-1.499));
    printf("Trunc (double): %d\n", trunc(-1.500));

    printf("Floor (double): %d\n", floor(1.499));
    printf("Floor (double): %d\n", floor(1.500));
    printf("Floor (double): %d\n", floor(-1.499));
    printf("Floor (double): %d\n", floor(-1.500));

    printf("Ceil (double): %d\n", ceil(1.499));
    printf("Ceil (double): %d\n", ceil(1.500));
    printf("Ceil (double): %d\n", ceil(-1.499));
    printf("Ceil (double): %d\n", ceil(-1.500));

    printf("Round (double): %d\n", round(1.499));
    printf("Round (double): %d\n", round(1.500));
    printf("Round (double): %d\n", round(-1.499));
    printf("Round (double): %d\n", round(-1.500));

    printf("Round to 0 places (double): %f\n", round(1.499, 0));
    printf("Round to 0 places (double): %f\n", round(1.500, 0));
    printf("Round to 0 places (double): %f\n", round(-1.499, 0));
    printf("Round to 0 places (double): %f\n", round(-1.500, 0));
    printf("Round to 1 place (double): %f\n", round(1.049, 1));
    printf("Round to 1 place (double): %f\n", round(1.050, 1));
    printf("Round to 1 place (double): %f\n", round(-1.049, 1));
    printf("Round to 1 place (double): %f\n", round(-1.050, 1));
    printf("Round to 3 place (double): %f\n", round(1.499, 3));
    printf("Round to 3 place (double): %f\n", round(1.500, 3));
    printf("Round to 3 place (double): %f\n", round(-1.499, 3));
    printf("Round to 3 place (double): %f\n", round(-1.500, 3));
    printf("Round to 4 place (double): %f\n", round(1.499, 4));
    printf("Round to 4 place (double): %f\n", round(1.500, 4));
    printf("Round to 4 place (double): %f\n", round(-1.499, 4));
    printf("Round to 4 place (double): %f\n", round(-1.500, 4));

    printf("Deg2Rad: %f\n", degToRad(420.0));
    printf("Deg2Rad: %f\n", degToRad(42.678));
    printf("Deg2Rad: %f\n", degToRad(321.453));

    printf("Rad2Deg: %f\n", radToDeg(1.0));
    printf("Rad2Deg: %f\n", radToDeg(0.0));
    printf("Rad2Deg: %f\n", radToDeg(1.234567));

    printf("Sin (double): %f\n", fct::sin(78.345));
    printf("Sin (int): %f\n", fct::sin(23));
    printf("Sin (short): %f\n", fct::sin(-68s));
    printf("Sin (long): %f\n", fct::sin(359l));

    printf("Cos (double): %f\n", fct::cos(78.345));
    printf("Cos (int): %f\n", fct::cos(23));
    printf("Cos (short): %f\n", fct::cos(-68s));
    printf("Cos (long): %f\n", fct::cos(359l));
}