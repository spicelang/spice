// Converts a double to an int
f<int> toInt(double input) {
    // ToDo: Implement
    return 0;
}

// Converts a double to a short
f<short> toInt(double input) {
    // ToDo: Implement
    return (short) 0;
}

// Converts a double to a long
f<long> toInt(double input) {
    // ToDo: Implement
    return (long) 0;
}

// Converts a double to a byte
f<byte> toByte(double input) {
    // ToDo: Implement
    result = (byte) 0;
}

// Converts a double to a string
f<string> toString(double input) {
    // ToDo: Implement
    return "";
}

// Converts a double to a boolean
f<bool> toBool(double input) {
    return input >= 0.5;
}