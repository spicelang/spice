type Struct struct {
    heap int* heapInt
}

f<int> main() {
    int a;
    printf("%d", a);
}