p unusedProcedure() {
    printf("Hello World!");
}

f<int> main() {}