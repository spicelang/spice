f<int> main() {
    int a = 1;
    int b = ++2;
    printf("Calculation result: %d", a + b);
}