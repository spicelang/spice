import "source1" as s1;

f<int> main() {
    dyn s = s1::Vector{1};
    printf("Result: %d\n", s.i);
}