/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/net/socket" as socket;

f<int> main() {
    socket.Socket s = socket.openServerSocket(8080s, 2);
    printf("Error code: %d", s.errorCode);
    //s.close();
}*/


ext<int> usleep(int);

f<int> main() {
    byte* t1;
    byte* t2;
    byte* t3;

    t1 = thread {
        printf("Thread 1 started: %p\n", t1);
        usleep(2000 * 1000);
        printf("Thread 1 finished\n");
    };

    t2 = thread {
        printf("Thread 2 started\n");
        printf("Tid 1: %p\n", t1);
        join(t1, t3);
        printf("Thread 2 finished\n");
    };

    t3 = thread {
        printf("Thread 3 started\n");
        usleep(3000 * 1000);
        printf("Thread 3 finished\n");
    };

    join(t1, t2, t3);
    printf("Program finished\n");
}