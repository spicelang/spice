f<int> main() {
    char* s = "abc";
    printf("%s\n", cast<char*>(s));
}