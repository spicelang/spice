import "std/os/syscall";

f<int> main() {
    string str = "Hello World!\n";
    syscallWrite(FileDescriptor::STDOUT, str);
}
