ext f<byte*> malloc(int);

f<int> test(string input) {
    return 12;
}

f<int> main() {
    f<int>(string) testFct = test;
    //int i = testFct();
    //printf("Result: %d", i);
}