/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.String s1 = str.String("Test string");
}*/

f<int> main() {
    assert 1 == 1;
    printf("Unreachable");
}