ext f<int> usleep(int);

f<int> main() {
    printf("Starting one thread ...\n");
    thread {
        usleep(500 * 1000);
        printf("Hello from the thread 1\n");
    }
    thread {
        usleep(200 * 1000);
        printf("Hello from the thread 2\n");
    }
    usleep(1000 * 1000);
    printf("Hello from original\n");
}