ext<int> mkdir(char*, int);

f<int> createDir(string pathStr, int mode) {
    char* path = pathStr;
    return mkdir(path, mode);
}