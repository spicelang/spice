f<int> main() {
    printf("Test", 3);
}