type Fruit enum {
    APPLE,
    BANANA,
    MANGO,
    ORANGE
}

f<int> main() {
    printf("Test: %d", Fruit.ORANGE);
}