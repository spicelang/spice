ext f<heap byte*> malloc(unsigned long);
ext f<heap byte*> malloc(unsigned long);

f<int> main() {}