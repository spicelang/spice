import "os-test2" as s1;

f<int> main() {
    Vector<int> v = Vector<int>{};
    v.setData(12);
    printf("Data: %d\n", v.data);
    v.setData(1);
    printf("Data: %d\n", v.data);
}