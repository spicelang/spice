f<int> main() {
    int value0 = 2;
    int[5] intArray = { value0, 7, 4 };
    intArray[2] = 11;
    intArray[0] = 3;
    printf("Item 0: %d, item 2: %d, item 4: %d", intArray[0], intArray[2], intArray[4]);
}
