import "std/data/map";

f<int> main() {
    Map<string, int> map;
    map["test"] = 1;
}