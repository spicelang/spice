import "test3" as s2;

p test() {
    printf("p: %f", s2.getDouble());
}