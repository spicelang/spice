// Mathematical constants
public const double E = 2.7182818284590452354;
public const double LOG2E = 1.4426950408889634074;
public const double LOG10E = 0.43429448190325182765;

public const double LN2 = 0.69314718055994530942;
public const double LN10 = 2.30258509299404568402;

public const double PI = 3.14159265358979323846;
public const double PI_2 = 1.57079632679489661923;
public const double PI_4 = 0.78539816339744830962;

public const double SQRT_2 = 1.41421356237309504880;
public const double SQRT_E = 1.64872127070012814685;
public const double SQRT_PI = 1.7724538509055160273;
public const double SQRT_PHI = 1.27201964951406896425;