// Imports
import "std/text/print";
import "std/os/cmd";
import "std/io/cli-parser";

/**
 * Representation of the various cli options
 */
public type CliOptions struct {
    public String mainSourceFile // e.g. main.spice
    public String targetTriple   // In format: <arch><sub>-<vendor>-<sys>-<abi>
    public String targetArch
    public String targetVendor
    public String targetOs
    public bool execute = false
    public bool isNativeTarget = true
    public String cacheDir
    public String outputDir      // Where the object files go. Should always be a temp directory
    public String outputPath     // Where the output binary goes.
    public unsigned short compileJobCount = 0 // O for auto
    public bool ignoreCache = false
    public bool printDebugOutput = false
    public bool dumpCST = false
    public bool dumpAST = false
    public bool dumpIR = false
    public bool dumpAssembly = false
    public bool dumpSymbolTables = false
    public bool disableAstOpt = false
    public short optLevel = 2s // -O0 = 0, -O1 = 1, -O2 = 2, -O3 = 3, -Os = 4, -Oz = 5
    public bool generateDebugInfo = false
    public bool disableVerifier = false
    public bool testMode = false
}

/**
 * Helper class to setup the cli interface and command line parser
 */
public type CliInterface struct {
    CliParser cliParser
    public CliOptions cliOptions
    public bool shouldCompile = false
    public bool shouldInstall = false
    public bool shouldExecute = false
}

public p CliInterface.createInterface() {
    this.cliParser = CliParser("Spice", "Spice programming language");
    this.cliParser.setFooter("Copyright (c) Marc Auberer 2021-2023");

    // Add version flag
    this.cliParser.setVersion("Spice version 0.14.3\nbuilt by: GitHub Actions\n\n(c) Marc Auberer 2021-2023");

    // Create sub-commands
    this.addBuildSubcommand();
    this.addRunSubcommand();
    this.addInstallSubcommand();
    this.addUninstallSubcommand();

    // ToDo: extend
}

/**
 * Validates if all necessary cli options were provided.
 *
 * @throws InvalidCliOptionsException if there were an invalid combination of cli options provided
 */
public p CliInterface.validate() {
    if ((this.cliOptions.targetArch.isEmpty() && this.cliOptions.targetVendor.isEmpty() && this.cliOptions.targetOs.isEmpty()) ||
        (!this.cliOptions.targetArch.isEmpty() && !this.cliOptions.targetVendor.isEmpty() && !this.cliOptions.targetOs.isEmpty())) {
        // ToDo: throw cli error
    }

    // Error out when opt level > 0 and debug info enabled
    if (this.cliOptions.optLevel > 0 && this.cliOptions.generateDebugInfo) {
        // ToDo: throw cli error
    }
}

/**
 * Initialize the cli options based on the input of the user
 */
public p CliInterface.enrich() {
    // Propagate target information
    if this.cliOptions.targetTriple.isEmpty() && this.cliOptions.targetArch.isEmpty() {
        // ToDo: Extend
    }

    // Dump AST, IR and symbol table if all debug output is enabled
    if this.cliOptions.printDebugOutput {
        this.cliOptions.dumpAST = true;
        this.cliOptions.dumpIR = true;
        this.cliOptions.dumpSymbolTables = true;
    }
}

/**
 * Add build subcommand to cli interface
 */
p CliInterface.addBuildSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.createSubcommand("build", "Builds your Spice program and emits an executable");
    subCmd.addAlias("b");

    addCompileSubcommandOptions(subCmd);

    // --target-triple
    Option& targetOption = subCmd.addOption("--target", this.cliOptions.targetTriple, "Target triple for the emitted executable (for cross-compiling)");
    targetOption.addAlias("--target-triple");
    targetOption.addAlias("-t");
    // --target-arch
    Option& targetArchOption = subCmd.addOption("--target-arch", this.cliOptions.targetArch, "Target arch for emitted executable (for cross-compiling)");
    // --target-vendor
    Option& targetVendorOption = subCmd.addOption("--target-vendor", this.cliOptions.targetVendor, "Target vendor for emitted executable (for cross-compiling)");
    // --target-os
    Option& targetOsOption = subCmd.addOption("--target-os", this.cliOptions.targetOs, "Target OS for emitted executable (for cross-compiling)");

    // --output
    Option& outputOption = subCmd.addOption("--output", this.cliOptions.outputPath, "Set the output file path");
    outputOption.addAlias("-o");
    // --debug-info
    Option& debugInfoOption = subCmd.addOption("--debug-info", this.cliOptions.generateDebugInfo, "Generate debug info");
    debugInfoOption.addAlias("-g");
    // --disable-verifier
    Option& disableVerifierOption = subCmd.addOption("--disable-verifier", this.cliOptions.disableVerifier, "Disable LLVM module and function verification");
}

/**
 * Add run subcommand to cli interface
 */
p CliInterface.addRunSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.createSubcommand("run", "Builds your Spice program and runs it immediately");
    subCmd.addAlias("r");

    addCompileSubcommandOptions(subCmd);

    // --output
    Option& outputOption = subCmd.addOption("--output", this.cliOptions.outputPath, "Set the output file path");
    outputOption.addAlias("-o");
    // --debug-info
    Option& debugInfoOption = subCmd.addOption("--debug-info", this.cliOptions.generateDebugInfo, "Generate debug info");
    debugInfoOption.addAlias("-g");
    // --disable-verifier
    Option& disableVerifierOption = subCmd.addOption("--disable-verifier", this.cliOptions.disableVerifier, "Disable LLVM module and function verification");
}

/**
 * Add install subcommand to cli interface
 */
p CliInterface.addInstallSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.createSubcommand("install", "Builds your Spice program and installs it to a directory in the PATH variable");
    subCmd.addAlias("i");

    addCompileSubcommandOptions(subCmd);
}

/**
 * Add uninstall subcommand to cli interface
 */
p CliInterface.addUninstallSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.createSubcommand("uninstall", "Builds your Spice program and runs it immediately");
    subCmd.addAlias("d");

    addCompileSubcommandOptions(subCmd);
}

p CliInterface.addCompileSubcommandOptions(CliSubcommand& subCmd) {

}

/**
 * Start the parsing process
 *
 * @param argc Argument count
 * @param argv Argument vector
 * @return Return code
 */
public f<int> CliInterface.parse(int argc, string[] argv) {
    return this.cliParser.parse(argc, argv);
}

/**
 * Executes the built executable
 */
p CliInterface.runBinary() {
    // Print status message
    if this.cliOptions.printDebugOutput {
        println("Running executable ...\n");
    }

    // Run executable
    execCmd(this.cliOptions.outputPath.getRaw());
}