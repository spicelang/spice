import "std/type/byte" as byteTy;

f<int> main() {
    // toDouble()
    double asDouble = byteTy.toDouble((byte) 15);
    assert asDouble == 15.0;

    // toInt()
    int asInt = byteTy.toInt((byte) 9);
    assert asInt == 9;

    // toShort()
    short asShort = byteTy.toShort((byte) 6);
    assert asShort == 6s;

    // toLong()
    long asLong = byteTy.toLong((byte) 63);
    assert asLong == 63l;

    // toString()
    //string asString = byteTy.toString((byte) 13);
    //assert asString == "13";

    // toBool()
    bool asBool1 = byteTy.toBool((byte) 1);
    assert asBool1 == true;
    bool asBool2 = byteTy.toBool((byte) 0);
    assert asBool2 == false;

    printf("All assertions succeeded");
}