f<int> testFunc(int input) {
    result = 1;
    if (input > 1) {
        printf("true");
        return 0;
    }
    printf("false");
}

f<int> main() {
    printf("Result: %d", testFunc(1));
}