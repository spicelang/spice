type DemoStruct struct {
    int i
    long l
    short s
    string str
}

f<int> main() {
    printf("%d\n", typeid(4));
    printf("%d\n", typeid<int>());

    DemoStruct s = DemoStruct{123, 56l, 12s, "String"};
    printf("%d\n", typeid<DemoStruct>());
    printf("%d\n", typeid(s));
}