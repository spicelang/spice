// Add generic type definitions
type T dyn;
type U int|short|long;

/**
 * The Iterable interface must be implemented in order to be handled as an iterator by Spice. For instance, all elements,
 * implementing the Iterable interface can be looped over by a standard foreach loop.
 */
public type Iterable<T> interface {
    f<bool> hasNext();
    f<T> next();
    f<T&> get();
}

/**
 * A BasicIterator in Spice is a commonly used data structure, which serves as a tool to loop over other iteratable
 * data structures
 */
public type NumberIterator<U> struct : Iterable<U> {
    U lowerBound
    U upperBound
    unsigned long index
}

public p NumberIterator.ctor(U lowerBound, U upperBound) {
    this.lowerBound = lowerBound;
    this.upperBound = upperBound;
    this.index = 0;
}

public inline const f<bool> NumberIterator.hasNext() {
    return this.lowerBound + this.index <= this.upperBound;
}

public inline f<U*> NumberIterator.next() {
    assert this.hasNext();
    this.index++;
    return this.data;
}

public inline f<U&> NumberIterator.get() {
    return this.lowerBound + this.index;
}