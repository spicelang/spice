// Std imports
import "std/data/unordered-map";

// Own imports

public type TypeRegistry struct {

}