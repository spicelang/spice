p test<byte>() {}

f<int> main() {
    test<int>();
}