p test(int param) {
    {
        {
            {
                {}
                printf("Param: %d\n", param);
                {}
            }
        }
    }
}

f<int> main() {
    test(12);
}