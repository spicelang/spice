type StructToCopy struct {
    heap int* intHeapPtr
}

f<int> main() {
    StructToCopy stc;
}
