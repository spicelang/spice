f<int> fib(int n) {
    if n <= 1 { return 1; }
    return fib(n - 1) + fib(n - 2);
}

f<int> main() {
    printf("Result: %d", fib(46));
}