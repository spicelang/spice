type Inner struct {
    short x = -43s
}

p Inner.ctor(const Inner& other) {
    this.x = other.x + 5s;
}

type Middle struct {
    Inner inner
}

type Outer struct {
    Middle middle
}

f<int> main() {
    Outer outer;
    printf("x = %d\n", outer.middle.inner.x);
    Outer outer2 = outer;
    printf("x = %d\n", outer2.middle.inner.x);
}