import "std/os/dir" as dir;

f<int> main() {
    //dir.mkDir("./test.txt");
}