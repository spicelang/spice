/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/net/socket" as socket;

f<int> main() {
    socket.Socket s = socket.openServerSocket(8080s, 2);
    printf("Error code: %d", s.errorCode);
    //s.close();
}*/

import "std/io/dir" as dir;

f<int> main() {
    printf("Existing before create: %d\n", dir.dirExists("./test"));
    dyn mkReturnCode = dir.mkDir("./test", dir.MODE_ALL_RWX);
    printf("mkDir return code: %d\n", mkReturnCode);
    printf("Existing after create: %d\n", dir.dirExists("./test"));
    dyn rmReturnCode = dir.rmDir("./test");
    printf("rmDir return code: %d\n", rmReturnCode);
    printf("Existing after delete: %d\n", dir.dirExists("./test"));
}