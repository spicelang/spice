// Std imports
import "std/data/unordered-map";

// Own imports
import "bootstrap/source-file-intf";
import "bootstrap/util/system-util";
import "bootstrap/global/global-resource-manager-intf";

// Constants
const string STRING_RT_IMPORT_NAME = "__rt_string";
const string RESULT_RT_IMPORT_NAME = "__rt_result";
const string ERROR_RT_IMPORT_NAME = "__rt_error";
const string MEMORY_RT_IMPORT_NAME = "__rt_memory";
const string RTTI_RT_IMPORT_NAME = "__rt_rtti";

public type RuntimeModule enum {
    STRING_RT = 1,
    RESULT_RT = 2,
    ERROR_RT  = 4,
    MEMORY_RT = 8,
    RTTI_RT   = 16
}

type ModuleNamePair struct {
    string importName
    string fileName
}

public type RuntimeModuleManager struct {
    IGlobalResourceManager &resourceManager
    UnorderedMap<RuntimeModule, ISourceFile *> modules
}

public p RuntimeModuleManager.ctor(IGlobalResourceManager &resourceManager) {
    this.resourceManager = resourceManager;
}

public f<ISourceFile *> RuntimeModuleManager.requestModule(ISourceFile* parentSourceFile, RuntimeModule requestedModule) {
    const String importName = String(this.resolveNamePair(requestedModule).importName);

    // Check if the requested module is available already, if not load it
    dyn rtFile = this.isModuleAvailable(requestedModule) ? this.getModule(requestedModule) : this.loadModule(parentSourceFile, requestedModule);

    // Add the dependency to the parent source file
    parentSourceFile.addDependency(rtFile, parentSourceFile.ast, importName, rtFile.filePath.toString());
    assert parentSourceFile.dependencies.contains(importName);
    ISourceFile* runtimeFile = parentSourceFile.dependencies.get(importName);
    this.modules.upsert(requestedModule, runtimeFile);

    // Merge the module name registry with the one of the source file
    parentSourceFile.mergeNameRegistries(*rtFile, importName);

    // Tell the source file, that the requested runtime has been imported
    parentSourceFile.importedRuntimeModules |= requestedModule;

    return runtimeFile;
}

public f<ISourceFile *> RuntimeModuleManager.getModule(RuntimeModule requestedModule) {
    assert this.modules.contains(requestedModule);
    return this.modules.get(requestedModule);
}

public f<bool> RuntimeModuleManager.isModuleAvailable(RuntimeModule requestedModule) {
    return this.modules.contains(requestedModule);
}

public f<ISourceFile *> RuntimeModuleManager.loadModule(ISourceFile* parentSourceFile, RuntimeModule requestedModule) {
    const ModuleNamePair namePair = this.resolveNamePair(requestedModule);
    const FilePath filePath = getStdDir() / "runtime" / namePair.fileName / ".spice";
    assert filePath != parentSourceFile.filePath;

    // Instruct the global resource manager to create a new source file
    SourceFile* moduleSourceFile = this.resourceManager.createSourceFile(parentSourceFile, namePair.importName, filePath, true);
    moduleSourceFile.isMainFile = false;

    // Run frontend and first type checker run for the loaded source file
    moduleSourceFile.runFrontEnd();
    moduleSourceFile.runTypeCheckerPre();

    return moduleSourceFile;
}

public f<ModuleNamePair> RuntimeModuleManager.resolveNamePair(RuntimeModule requestedModule) {
    switch requestedModule {
        case RuntimeModule::STRING_RT: {
            return ModuleNamePair{STRING_RT_IMPORT_NAME, "string_rt"};
        }
        case RuntimeModule::RESULT_RT: {
            return ModuleNamePair{RESULT_RT_IMPORT_NAME, "result_rt"};
        }
        case RuntimeModule::ERROR_RT: {
            return ModuleNamePair{ERROR_RT_IMPORT_NAME, "error_rt"};
        }
        case RuntimeModule::MEMORY_RT: {
            return ModuleNamePair{MEMORY_RT_IMPORT_NAME, "memory_rt"};
        }
        case RuntimeModule::RTTI_RT: {
            return ModuleNamePair{RTTI_RT_IMPORT_NAME, "rtti_rt"};
        }
        default: {
            panic(Error("Requested unknown runtime module"));
        }
    }
}