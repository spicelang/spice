type TestStruct struct {
    double dbl
    string* str
    bool bl
}

f<int> main() {
    dyn str = "Hello!";
    dyn testInstance = TestStruct { &str, false };
    printf("Double: %f", testInstance.dbl);
}