// Link external functions
ext f<heap byte*> malloc(long);
ext p free(heap byte*);

// Add generic type definitions
type T dyn;

/**
 * Node of a LinkedList
 */
public type Node<T> struct {
    T value
    heap Node<T>* next
}

/**
 * A linked list is a common, dynamically resizable data structure to store uniform data in order.
 * It is characterized by the pointer for each item, pointing to the next one.
 *
 * E.g. for a LinkedList<int>:
 * 1234 -> 4567 -> 7890 -> 4567 -> nil<int*>
 * tail                    head
 *
 * Time complexity:
 * Insert: O(1)
 * Delete: O(1)
 * Search: O(n)
 *
 * Beware that each add operation allocates memory and every remove operation frees memory.
 */
public type LinkedList<T> struct {
    heap Node<T>* tail
    heap Node<T>* head
}

public p LinkedList.ctor() {
    this.tail = nil<heap Node<T>*>;
    this.head = nil<heap Node<T>*>;
}

public p LinkedList.dtor() {
    Node<T>* curr = this.tail;
    while curr != nil<heap Node<T>*> {
        Node<T>* next = curr.next;
        free(curr);
        curr = next;
    }
}

public p LinkedList.insert(const T& value) {
    // Create new node
    heap Node<T>* newNode;
    unsafe {
        newNode = (heap Node<T>*) malloc(sizeof(type Node<T>) / 8l);
    }
    newNode.value = value;
    newNode.next = nil<heap Node<T>*>;

    // Insert at head
    this.head.next = newNode;
    this.head = newNode;
}

public p LinkedList.insertAt(unsigned long idx, const T& value) {
    // Create new node
    heap Node<T>* newNode;
    unsafe {
        newNode = (heap Node<T>*) malloc(sizeof(type Node<T>) / 8);
    }
    newNode.value = value;

    // Search for item right before insert position
    Node<T>* prev = this.tail;
    while curr != nil<heap Node<T>*> && idx > 1 {
        prev = prev.next;
        idx--;
    }

    // Link the next node to the new one
    newNode.next = prev.next;
    // Link the new node to the previous one
    prev.next = newNode;

    // Check if we have a new tail
    if idx == 0l {
        this.tail = newNode;
    }
    // Check if the previous node was the last node
    if this.head == prev {
        this.head = newNode;
    }
}

public p LinkedList.remove(const T& valueToRemove) {
    heap Node<T>* curr = this.tail;
    heap Node<T>* prev = nil<heap T*>;
    while curr != nil<heap Node<T>*> && curr.value != valueToRemove {
        prev = curr;
        curr = curr.next;
    }
    // Check if the item was found. If yes, delete its node
    if curr != nil<heap Node<T>*> {
        // Set the next node of the previous node
        prev.next = curr.next;
        // Free the removed node
        free(curr);
    }
}

public inline f<T&> LinkedList.getFirst() {
    return this.head.value;
}

public inline f<T&> LinkedList.getLast() {
    return this.tail.value;
}