type TestStruct struct {
    unsigned int field1
    long field2
}

f<int> main() {
    printf("Size: %d\n", sizeof(TestStruct{}));
}