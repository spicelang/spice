/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec.Vector<pair.Pair<int, string>> pairVector = vec.Vector<pair.Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair.Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

p testProc(int[]*** nums) {
    int[]* nums1 = **nums;
    int[] nums2 = *nums1;
    nums2[2] = 10;
    printf("1: %d\n", nums2[0]);
    printf("2: %d\n", nums2[1]);
    printf("3: %d\n", nums2[2]);
    printf("4: %d\n", nums2[3]);
}

f<int> main() {
    int[4] intArray = { 1, 2, 3, 4 };
    printf("1: %d\n", intArray[1]);
    testProc(&&&intArray);
}