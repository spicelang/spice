ext<dyn> exteralFunction();

f<int> main() {
    externalFunction(1, 3);
}