import "std/data/unordered-map";

f<int> main() {
    UnorderedMap<int, string> map;
    map.upsert(1, "one");
    map.upsert(2, "two");
    map.upsert(3, "three");
    assert map.contains(1);
    assert map.contains(2);
    assert map.contains(3);
    assert !map.contains(4);
    assert map.getSize() == 3;
    for int i = 1; i <= 3; i++ {
        printf("%s\n", map.get(i));
    }
    const Result<string> item4 = map.getSafe(4);
    assert item4.isErr();
    map.remove(2);
    assert !map.contains(2);
    assert map.getSize() == 2;
    map.clear();
    assert map.getSize() == 0;


    printf("All assertions passed!\n");
}

/*import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

f<int> main() {
    DefaultMemoryManager defaultMemoryManager;
    IMemoryManager* memoryManager = &defaultMemoryManager;
    BlockAllocator<int> allocator = BlockAllocator<int>(memoryManager, 10l);
}*/