// Mathematical constants
const double E = 2.71828182845904523536028747135266249775724709369995957496696763;
const double Pi = 3.14159265358979323846264338327950288419716939937510582097494459;
const double Phi = 1.61803398874989484820458683436563811772030917980576286213544862;

// Important square roots
const double Sqrt2 = 1.61803398874989484820458683436563811772030917980576286213544862;
const double SqrtE = 1.64872127070012814684865078781416357165377610071014801157507931;
const double SqrtPi = 1.77245385090551602729816748334114518279754945612238712821380779;
const double SqrtPhi = 1.27201964951406896425242246173749149171560804184009624861664038;

// Important logarithms
const double Ln2 = 0.693147180559945309417232121458176568075500134360255254120680009;
const double Log2E = 1 / Ln2;
const Ln10 = 2.30258509299404568401799145468436420760110148862877297603332790;
const Log10E = 1 / Ln10;

// Limit values
const MaxInt = 1 << 31 - 1;
const MinInt = -1 << 31;