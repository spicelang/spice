//import "std/type/int" as unused;
//import "os-test2" as s1;

type TestStruct struct {
    int field1
    double field2
}

p TestStruct.ctor() {
    this.field1 = 1;
}

f<int> main() {
    dyn testStruct = TestStruct(345);
}