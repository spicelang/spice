// Constants
const unsigned long INITIAL_ALLOC_COUNT = 5l;
const unsigned int RESIZE_FACTOR = 2;

// Link external functions
ext<byte*> malloc(long);
ext<byte*> realloc(byte*, int);
ext free(byte*);
ext<byte*> memcpy(byte*, byte*, int);

// Add generic type definition
type T dyn;

/**
 * A queue in Spice is a commonly used data structure, which uses the FiFo (first in, first out) principle
 */
public type Queue<T> struct {
    T* contents             // Pointer to the first data element
    unsigned long capacity  // Allocated number of items
    unsigned long size      // Current number of items
    unsigned long idxFront  // Index for front access
    unsigned long idxBack   // Index for back access
    unsigned int itemSize   // Size of a single item
}

public p Queue.ctor(unsigned long initAllocItems, const T& defaultValue) {
    // Allocate space for the initial number of elements
    this.ctor(initAllocItems);
    // Fill in the default values
    for int index = 0; index < initAllocItems; index++ {
        unsafe {
            this.contents[index] = defaultValue;
        }
    }
    this.size = initAllocItems;

}

public p Queue.ctor(unsigned int initAllocItems) {
    this.ctor((long) initAllocItems);
}

public p Queue.ctor(unsigned long initAllocItems = INITIAL_ALLOC_COUNT) {
    // Allocate space for the initial number of elements
    this.itemSize = sizeof(type T) / 8;
    unsafe {
        this.contents = (T*) malloc(this.itemSize * initAllocItems);
    }
    this.size = 0l;
    this.capacity = initAllocItems;
    this.idxFront = 0l;
    this.idxBack = 0l;
}

public p Queue.dtor() {
    // Free all the memory
    unsafe {
        free((byte*) this.contents);
    }
}

/**
 * Add an item at the end of the queue
 */
public p Queue.push(const T& item) {
    // Check if we need to re-allocate memory
    if this.isFull() {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Insert the element at the back
    unsafe {
        this.contents[(int) this.idxBack++] = item;
    }

    // Increase size
    this.size++;
}

/**
 * Retrieve the first item and remove it
 *
 * @return First item
 */
public f<T&> Queue.pop() {
    this.size--;
    unsafe {
        return this.contents[(int) this.idxFront++];
    }
}

/**
 * Retrieve the first item without removing it from the queue
 *
 * @return First item
 */
public f<T&> Queue.front() {
    assert !this.isEmpty();
    unsafe {
        return this.contents[(int) this.idxFront];
    }
}

/**
 * Retrieve the last item without removing it from the queue
 *
 * @return Last item
 */
public f<T&> Queue.back() {
    assert !this.isEmpty();
    unsafe {
        return this.contents[(int) this.idxBack];
    }
}

/**
 * Retrieve the current size of the queue
 *
 * @return Current size of the queue
 */
public f<long> Queue.getSize() {
    return this.size;
}

/**
 * Retrieve the current capacity of the queue
 *
 * @return Current capacity of the queue
 */
 public f<long> Queue.getCapacity() {
     return this.capacity;
 }

/**
 * Checks if the queue contains any items at the moment
 *
 * @return Empty or not empty
 */
public f<bool> Queue.isEmpty() {
    return this.size == 0;
}

/**
 * Checks if the queue exhausts its capacity and needs to resize at the next call of push
 *
 * @return Full or not full
 */
public f<bool> Queue.isFull() {
    return this.size == this.capacity;
}

/**
 * Reserves `itemCount` items
 */
public p Queue.reserve(unsigned long itemCount) {
    if itemCount > this.capacity {
        this.resize(itemCount);
    }
}

/**
 * Frees allocated memory that is not used by the queue
 */
public p Queue.pack() {
    // Return if no packing is required
    if this.isFull() { return; }
    // Pack the array
    this.resize(this.size);
}

/**
 * Re-allocates heap space for the queue contents
 */
p Queue.resize(unsigned long itemCount) {
    // Allocate the new memory
    unsafe {
        byte* oldAddress = (byte*) this.contents;
        int newSize = (int) (this.itemSize * itemCount);
        T* newMemory = (T*) realloc(oldAddress, newSize);
        this.contents = newMemory;
    }
    // Set new capacity
    this.capacity = itemCount;
}