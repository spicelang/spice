/**
 * Asserts that a condition evaluates to true. If that is not the case, the program will terminate with the passed error message
 *
 * @param condition Condition to check
 * @param message Message to print if the condition evaluates to false
 */
public p assertCondition(bool condition, string message = "<no-message>") {
    if (!condition) {

    }
}

/**
 * Concatenate two strings and return the concatenated result
 *
 * @param a part 1 of the result
 * @param b part 2 of the result
 *
 * @return Concatenated string
 */
public f<string> concat(string a, string b) {
    // Get wrapped instances of the raw strings
    String aWrapped = String(a);
    String bWrapped = String(b);
    // Append b to a
    aWrapped.append(bWrapped);
    // Return the raw outcome
    return aWrapped.getRaw();
}