import "source" as s;

p test() {
    printf("p: %f", s.getDouble());
}