f<int> main() {
    int[10] intArray = { 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 };
    foreach int i = 3, int item : intArray {
        printf("Array item no. %d: %d, ", i, item);
        i += 2;
    }
}