f<dyn> test() {
    return 1;
}

f<int> main() {
    dyn t = test();
}