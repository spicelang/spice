/*f<int> main() {
    int value0 = 2;
    int[5] intArray = { value0, 7, 4 };
    intArray[2] = 11;
    intArray[0] = 3;
    printf("Array item 0: %d, array item 2: %d", intArray[0], intArray[2]);
}*/

f<int> main() {
    string food = "Pizza";
    string* ptr = &food;

    printf("Pointer address: %p, value: %s", ptr, *ptr);

    /*ptr = "Burger";

    dyn restoredFood = *ptr;
    printf("Restored value: %s", restoredFood);

    printf("Restored value address: %p", &restoredFood);*/
}