import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = new str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();

    /*string a = "Hello";
    string b = "World";

    string c = a + " " + b + "!";
    printf("Concatenated string: %s\n", c);*/
}