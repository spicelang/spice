f<int> fibo(int n) {
    if n <=1 {
        return n;
    }
    return fibo(n-1) + fibo(n-2);
}

f<int> main() {
    sout.print(fibo(5));
}