f<int> main() {
    int test = 12;
    int* testPtr = &test;
    int test1 = testPtr;
    printf("Value1: %d, pointer: %p, value: %d", test, testPtr, test1);
}