// Imports
import "std/text/analysis";
import "std/math/fct";
import "std/type/type-conversion";

// Constants
const unsigned int ASCII_SHIFT_OFFSET = 32;
const char MIN_LOWER_CHAR = 'a';
const char MAX_LOWER_CHAR = 'z';
const char MIN_UPPER_CHAR = 'A';
const char MAX_UPPER_CHAR = 'Z';

// Generic type defs
type IntLongShort int|long|short;

/**
 * Returns the given char as upper case version
 *
 * @return Char in upper case
 */
public f<char> toUpper(char c) {
    if c >= MIN_LOWER_CHAR && c <= MAX_LOWER_CHAR {
        c -= cast<char>(ASCII_SHIFT_OFFSET);
    }
    return c;
}

/**
 * Returns the given text in caps
 *
 * @return Text in caps
 */
public f<String> toUpper(const String& text) {
    result = text;
    for unsigned long i = 0l; i < result.getLength(); i++ {
        result[i] = toUpper(result[i]);
    }
}

/**
 * Returns the given char as lower case version
 *
 * @return Char in lower case
 */
public f<char> toLower(char c) {
    if c >= MIN_UPPER_CHAR && c <= MAX_UPPER_CHAR {
        c += cast<char>(ASCII_SHIFT_OFFSET);
    }
    return c;
}

/**
 * Returns the given text in all-lower letters
 *
 * @return Text in all-lower letters
 */
public f<String> toLower(const String& text) {
    result = text;
    for unsigned long i = 0l; i < result.getLength(); i++ {
        result[i] = toLower(result[i]);
    }
}

/**
 * Returns the given text in capitalized form
 *
 * @return Capitalized text
 */
public f<String> capitalize(const String& text) {
    result = text;
    if result.getLength() >= 1 {
        result[0] = toUpper(result[0]);
    }
}

/**
 * Format the given number with thousands delimiter
 *
 * @param input Number
 * @param delimiter Custom thousands delimiter
 * @return Formatted string
 */
public f<String> formatThousandsDelimiter(int input, char delimiter = ',') {
    result = toString(input);
    const unsigned long n = result.getLength();
    const bool isNegative = input < 0;

    long insertPosition = n - 3;
    long stopPosition = isNegative ? 1l : 0l;
    while insertPosition > stopPosition {
        result.insert(insertPosition, delimiter);
        insertPosition -= 3;
    }
}

/**
 * Returns a formatted storage string (e.g. 1.4 MB for 1,500,000)
 *
 * @param bytes Number of bytes
 * @param useFactor1024 Use factor 1024 instead the default factor of 1000
 * @return Formatted string
 */
public f<String> formatStorageSize(unsigned long bytes, bool useFactor1024 = false) {
    const string[7] storageUnits1000 = ["B", "KB",  "MB",  "GB",  "TB",  "PB",  "EB"];
    const string[7] storageUnits1024 = ["B", "KiB", "MiB", "GiB", "TiB", "PiB", "EiB"];
    assert len(storageUnits1000) == len(storageUnits1024); // Sanity check

    const string[7]& storageUnits = useFactor1024 ? storageUnits1024 : storageUnits1000;
    const unsigned int factor = useFactor1024 ? 1024 : 1000;

    double size = cast<double>(bytes);
    unsigned int unitIndex = 0u;
    while size >= factor && unitIndex < len(storageUnits1000) {
        size /= cast<double>(factor);
        unitIndex++;
    }

    const double sizeRounded = round(size, 2);
    return toString(sizeRounded) + ' ' + storageUnits[unitIndex];
}
