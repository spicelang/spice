import "std/type/string" as str;

// Constants
const unsigned long INITIAL_ALLOC_COUNT = 5l;
const unsigned int RESIZE_FACTOR = 2;

// Link external functions
ext<byte*> malloc(long);
ext<byte*> realloc(byte*, int);
ext free(byte*);
ext<byte*> memcpy(byte*, byte*, int);

/**
 * String wrapper for enriching raw strings with information and make them mutable
 */
public type String struct {
    char* contents   // Pointer to the first char
    unsigned long capacity     // Allocated number of chars
    unsigned long length       // Current number of chars
}

public p String.ctor(string value = "") {
    // Allocate space for the initial number of elements
    int itemSize = sizeof(type char);
    unsafe {
        this.contents = (char*) malloc(itemSize * INITIAL_ALLOC_COUNT);
    }
    this.length = str.getRawLength(value);
    this.capacity = INITIAL_ALLOC_COUNT;
}

public p String.dtor() {
    // Free all the memory
    unsafe {
        free((byte*) this.contents);
    }
}

/**
 * Appends the given string wrapper to the current one
 *
 * @param appendix String wrapper to be appended
 */
public p String.append(String appendix) {
    for int i = 0; i < appendix.length; i++ {
        char charToAppend;
        unsafe {
            charToAppend = appendix.contents[i];
        }
        this.appendChar(charToAppend);
    }
}

/**
 * Appends the given char to the string and resize it if needed
 *
 * @param c Char to append
 */
public p String.appendChar(char c) {
    // Check if we need to re-allocate memory
    if this.length == this.capacity {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Insert the char at the right position
    unsafe {
        this.contents[this.length++] = c;
    }
}

/**
 * Get the raw and immutable string from this container instance
 *
 * @return Raw immutable string
 */
public f<string> String.getRaw() {
    return (string) this.contents;
}

/**
 * Retrieve the current length of the string
 *
 * @return Current length of the string
 */
public f<long> String.getLength() {
    return this.length;
}

/**
 * Retrieve the current capacity of the string
 *
 * @return Current capacity of the string
 */
 public f<long> String.getCapacity() {
     return this.capacity;
 }

/**
 * Checks if the string exhausts its capacity
 *
 * @return Full or not full
 */
public f<bool> String.isFull() {
    return this.length == this.capacity;
}

/**
 * Replaces the current contents of the string with an empty string
 */
public p String.clear() {
    this.length = 0l;
}

/**
 * Reserves `charCount` items
 */
public p String.reserve(unsigned long charCount) {
    if charCount > this.capacity {
        this.resize(charCount);
    }
}

/**
 * Re-allocates heap space for the string contents
 *
 * @param newLength new length of the string after resizing
 */
p String.resize(unsigned long newLength) {
    // Allocate the new memory
    unsafe {
        byte* oldAddress = (byte*) this.contents;
        int newSize = (int) (sizeof(type char) * newLength);
        char* newMemory = (char*) realloc(oldAddress, newSize);
        this.contents = newMemory;
    }
    // Set new capacity
    this.capacity = newLength;
}