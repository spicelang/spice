type Size alias unsigned long;