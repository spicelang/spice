f<int> testFunction(int arg0, dyn arg1 = "value", dyn arg2) {
    return 1;
}

f<int> main() {
    testFunction(12345);
}