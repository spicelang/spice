f<int> testFunc() {
    printf("Test func 1\n");
    return 1;
}

f<int> testFunc(string param) {
    printf("Test func 2: %s\n", param);
    return 2;
}

f<int> main() {
    int res = testFunc();
    printf("Result: %d\n", res);
    res = testFunc("param value");
}