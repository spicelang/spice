public const int SIZE = 16;
public const short MIN_VALUE = -32768s;
public const short MAX_VALUE = 32767s;

// External functions
ext f<unsigned int> snprintf(char*, unsigned long, string, short);

// Converts a short to a double
public f<double> toDouble(short input) {
    return 0.0 + input;
}

// Converts a short to an int
public f<int> toInt(short input) {
    return (int) input;
}

// Converts a short to a long
public f<long> toLong(short input) {
    return (long) input;
}

// Converts a short to a byte
public f<byte> toByte(short input) {
    return (byte) ((int) input);
}

// Converts a short to a char
public f<char> toChar(short input) {
    return (char) input;
}

// Converts a short to a string
public f<String> toString(short input) {
    const unsigned int length = snprintf(nil<char*>, 0l, "%hd", input);
    result = String(length);
    snprintf((char*) result.getRaw(), length + 1l, "%hd", input);
}

// Converts a short to a boolean
public f<bool> toBool(short input) {
    return input >= 1;
}

// Check if the input is a power of two
public f<bool> isPowerOfTwo(short input) {
    return (input & (input - 1s)) == 0s;
}