f<int> main() {
    int test = 123;
    int& testRef = test;
    assert &test == &testRef;
}

/*ext<byte*> malloc(long);
ext free(byte*);

f<int> main() {
    byte* address = malloc(1l);
    *address = (byte) 12;
    free(address);
}*/

/*f<int> main() {
    int[10] a;
    for int i = 0; i < len(a); i++ {
        a[i] = 1;
    }
    printf("Cell [3]: %d", a[3]);
}*/