type UnusedStruct struct {
    double f1
    int* f2
}

f<int> main() {
    printf("%p", UnusedStruct{}.f2);
}