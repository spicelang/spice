f<int> main() {
    long alignment = alignof(type Test);
    printf("Alignment: %d", alignment);
}