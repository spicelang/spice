import "std/iterators/iterable";
import "std/data/vector";

// Generic type definitions
type T dyn;

/**
 * Iterator to iterate over a vector data structure
 */
public type VectorIterator<T> struct : Iterable<T> {
    Vector<T>& vector
    unsigned long cursor
}

public p VectorIterator.ctor<T>(Vector<V>& vector) {
    this.vector = vector;
    this.cursor = 0l;
}

/**
 * Check if the vector has another item
 *
 * @return true or false
 */
public inline const f<bool> VectorIterator.hasNext() {
    return this.cursor < this.vector.getSize();
}

/**
 * Returns the current item of the vector iterator and moves the cursor to the next item
 *
 * @return current item
 */
public inline f<T&> VectorIterator.next() {
    assert this.hasNext();
    T currentItem = this.get();
    this.cursor++;
    return currentItem;
}

/**
 * Returns the current item of the vector iterator
 */
public inline f<T&> VectorIterator.get() {
    return this.vector.get(this.cursor);
}