type T int|long|short;

type CompareResult enum {
    LESS,
    EQUAL,
    GREATER
}

type Compareable<T> interface {
    f<CompareResult> compare<T>(const T&, const T&);
}

type Person struct : Compareable<long> {
    string _firstName
    string _lastName
    unsigned int _age
}

f<CompareResult> Person.compare(const long& a, const long& b) {
    if a > b { return CompareResult::GREATER; }
    if a < b { return CompareResult::LESS; }
    return CompareResult::EQUAL;
}

f<int> main() {
    Person mike = Person{ "Mike", "Miller", 43 };
    const bool isEqual = mike.compare(22l, 22l) == CompareResult::EQUAL;
    printf("%d", isEqual);
}