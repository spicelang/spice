// Std imports

// Own imports

public type ISourceFile interface {

}