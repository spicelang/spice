type TestStruct struct {
    int* field1
    double field2
}

f<int> main() {
    int input = 12;
    dyn instance = new TestStruct { &input, 46.34 };
    TestStruct instance1 = instance;
    printf("Field1: %p, field2: %f", instance1.field1, instance1.field2);
}