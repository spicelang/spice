import "std/test/lifetime-object";

f<LifetimeObject> spawnLO() {
    return LifetimeObject();
}

f<int> main() {
    // Ignored return value of ctor
    printf("Ignored return value of ctor:\n");
    {
        LifetimeObject();
    }

    // Normal lifecycle
    printf("Normal lifecycle:\n");
    {
        LifetimeObject lo = LifetimeObject(); // ctor call
        LifetimeObject loCopy = lo; // copy ctor call
    } // dtor calls for both lo and loCopy at end of scope

    // Return from lambda as value
    printf("Return from lambda as value:\n");
    {
        const f<LifetimeObject>() spawnLO = f<LifetimeObject>() {
            return LifetimeObject();
        };

        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    // Return from lambda as reference
    printf("Return from lambda as reference:\n");
    {
        LifetimeObject loOrig = LifetimeObject();
        const f<LifetimeObject&>() spawnLO = f<LifetimeObject&>() {
            return loOrig;
        };

        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    // Return from lambda as const reference
    printf("Return from lambda as const reference:\n");
    {
        LifetimeObject loOrig = LifetimeObject();
        const f<const LifetimeObject&>() spawnLO = f<const LifetimeObject&>() {
            return loOrig;
        };

        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    // Return from function as value
    printf("Return from function as value:\n");
    {
        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    printf("Ternary (true temporary, false temporary)\n");
    {
        bool cond = true;
        LifetimeObject loCopy1 = cond ? LifetimeObject() : LifetimeObject(); // ctor calls in both branches
        LifetimeObject loCopy2 = !cond ? LifetimeObject() : LifetimeObject(); // ctor calls in both branches
    }

    printf("Ternary (true temporary, false not temporary)\n");
    {
        bool cond = true;
        LifetimeObject lo = LifetimeObject();
        LifetimeObject loCopy1 = cond ? LifetimeObject() : lo; // ctor in true branch, copy ctor in false branch
        LifetimeObject loCopy2 = !cond ? LifetimeObject() : lo; // ctor in true branch, copy ctor in false branch
    }

    printf("Ternary (true not temporary, false temporary)\n");
    {
        bool cond = true;
        LifetimeObject lo = LifetimeObject();
        LifetimeObject loCopy1 = cond ? lo : LifetimeObject(); // copy ctor in true branch, ctor in false branch
        LifetimeObject loCopy2 = !cond ? lo : LifetimeObject(); // copy ctor in true branch, ctor in false branch
    }

    printf("Ternary (true not temporary, false not temporary)\n");
    {
        bool cond = true;
        LifetimeObject lo1 = LifetimeObject();
        LifetimeObject lo2 = LifetimeObject();
        LifetimeObject loCopy1 = cond ? lo1 : lo2; // copy ctor call in both branches
        LifetimeObject loCopy2 = !cond ? lo1 : lo2; // copy ctor call in both branches
    }
}