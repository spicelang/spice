f<int> main() {
    double loopCounterOuter = 0.0;
    while (loopCounterOuter < 10) {
        loopCounterOuter += 0.15;
        if (loopCounterOuter < 4) {
            short loopCounterInner = 10s;
            while (loopCounterInner > 0) {
                printf("Outer: %f, inner: %d\n", loopCounterOuter, loopCounterInner);
                loopCounterInner--;
                if (loopCounterInner == 5) {
                    continue 2;
                }
            }
        }
    }
}