// Generic type defs
type TT int|long|short|bool; // Trivially hashable types
type TC byte|char; // Trivially hashable types with one additional cast
type T dyn; // Any type

// Aliases
public type Hash alias unsigned long;

public type IHashable interface {
    public f<Hash> hash();
}

/**
 * Hash primitive numeric type
 *
 * @param input Primitieve numeric to hash
 * @return Hash of primitive numeric
 */
public f<Hash> hash<TT>(TT input) {
    return cast<Hash>(input);
}

/**
 * Hash primitive numeric type
 *
 * @param input Primitieve numeric to hash
 * @return Hash of primitive numeric
 */
public f<Hash> hash<TC>(TC input) {
    return cast<Hash>(cast<unsigned int>(input));
}

/**
 * Hash a double value
 *
 * @param input Double to hash
 * @return Hash of double
 */
public f<Hash> hash(double input) {
    unsafe {
        return *(cast<Hash*>(&input));
    }
}

/**
 * Hash contents of an immutable string
 *
 * @param input String to hash
 * @return Hash of string
 */
public f<Hash> hash(string input) {
    // Hash using djb2 algorithm
    Hash hash = 5381l;
    for unsigned long i = 0l; i < len(input); i++ {
        Hash c = cast<Hash>(cast<unsigned int>(input[i]));
        hash = ((hash << 5l) + hash) + c; // hash * 33 + c
    }
    return hash;
}

/**
 * Hash contents of a mutable String object
 *
 * @param input String to hash
 * @return Hash of string
 */
public f<Hash> hash(const String& input) {
    return hash(input.getRaw());
}

/**
 * Dispatch function for structs, that implement the IHashable interface
 *
 * @param hashable Hashable object
 * @return Hash of the struct
 */
public f<Hash> hash(const IHashable& hashable) {
    return hashable.hash();
}
