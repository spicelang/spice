public const int SIZE = 16;
public const short MIN_VALUE = -32768;
public const short MAX_VALUE = 32767;

// Converts a short to a double
public f<double> toDouble(short input) {
    return 0.0 + input;
}

// Converts a short to an int
public f<int> toInt(short input) {
    return (int) input;
}

// Converts a short to a long
public f<long> toLong(short input) {
    return (long) input;
}

// Converts a short to a byte
public f<byte> toByte(short input) {
    return (byte) input;
}

// Converts a short to a char
public f<char> toChar(short input) {
    return (char) input;
}

// Converts a short to a string
public f<string> toString(short input) {
    // ToDo: Implement (See https://github.com/golang/go/blob/master/src/strconv/itoa.go)
    return "";
}

// Converts a v to a boolean
public f<bool> toBool(v input) {
    return input >= 1;
}