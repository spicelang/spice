f<int> main() {
    switch 1 {
        case false: { return 1; }
        default: { return 0; }
    }
}
