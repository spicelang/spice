import "std/os/mutex";

// Generic type defs
type T dyn;

public type Atomic<T> struct {
    T value
    Mutex mutex
}

public p Atomic.ctor() {
    this.value = cast<T>(0);
}

public p Atomic.ctor(T value) {
    this.value = value;
}

public p Atomic.store(const T& value) {
    LockGuard _ = LockGuard(this.mutex);
    this.value = value;
}

public const f<const T&> Atomic.load() {
    LockGuard _ = LockGuard(this.mutex);
    return this.value;
}

public f<T> Atomic.exchange(const T& value) {
    LockGuard _ = LockGuard(this.mutex);
    T old = this.value;
    this.value = value;
    return old;
}

public f<bool> Atomic.compareExchange(const T& expected, const T& desired) {
    LockGuard _ = LockGuard(this.mutex);
    result = this.value == expected;
    if result {
        this.value = desired;
    }
}