type T int|double|short|long;

f<int> sumNumbers<T>(T[] numberArray, int arrayLength) {
    result = 0;
    for int i = 0; i < arrayLength; i++ {
        result += numberArray[i];
    }
}

f<int> main() {
    short[7] numberList1 = { 1s, 2s, 3s, 4s, 5s, 6s, 7s };
    int result1 = sumNumbers<short>(numberList1, sizeof(numberList1));

    long[4] numberList2 = { 10l, 12l, 14l, 16l };
    int result2 = sumNumbers<long,short>(numberList2, sizeof(numberList2));

    printf("Results: %d, %d\n", result1, result2);
}