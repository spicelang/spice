f<int> main() {
    printf("This is a double: %f", 5.6);
    printf("This is an int: %d", 5);
    dyn variable = "test";
    printf("This is a pointer: %p", &variable);
    printf("This is a string: %c", "test");
}