ext f<byte*> malloc(long);
ext p free(byte*);

f<int> main() {
    byte* address = malloc(1l);
    *address = cast<byte>(12);
    free(address);
}