#![core.linker.flag]

f<int> main() {}