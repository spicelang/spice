// Std imports
import "bootstrap/data/unordered-map";

// Own imports

public type TypeRegistry struct {

}