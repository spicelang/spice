f<int> main() {
    printf("Result: %d", sizeof(type int));
}