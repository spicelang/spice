import "std/iterators/ranges";

f<int> main() {
    foreach int i : range(1, 5) {
        printf("%d\n", i);
    }
    /*int i;
    for (dyn it = range(1, 5); it.hasNext(); i = it.next()) {
        printf("%d\n", i);
    }*/
}