f<int> main() {
    int& i = 123;
    printf("Hello: %d\n", i);
}