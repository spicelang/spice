/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec.Vector<pair.Pair<int, string>> pairVector = vec.Vector<pair.Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair.Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

ext<int> usleep(int);

f<int> main() {
    byte* t1;
    byte* t2;
    byte* t3;

    t1 = thread {
        usleep(300 * 1000);
        printf("Thread 1 finished\n");
    };

    t2 = thread {
        join(t1, t3);
        printf("Thread 2 finished\n");
    };

    t3 = thread {
        usleep(200 * 1000);
        printf("Thread 3 finished\n");
    };

    join(t1, t2, t3);
    printf("Program finished\n");
}