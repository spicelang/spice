f<string> testFunction() {
    return 7;
}

f<int> main() {
    testFunction();
    return 0;
}