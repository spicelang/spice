public type Driveable interface {
    public p drive(int);
    public f<bool> isDriving();
}