/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "socket" as socket;

f<int> main() {
    socket.Socket s = socket.openServerSocket(8080s);
    //socket.NestedSocket n = s.nested;
    //printf("%s", n.testString);
}*/


type TestStruct struct {
    string test
    int test1
}

f<int> TestStruct.compute() {
    string test = "Test";
    return this.test1;
}

f<int> main() {
    printf("%d", TestStruct{ "sdf", 12 }.compute());
}