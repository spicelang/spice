import "test" as test;