f<string> unusedReturnValue() {
    return "unused";
}

f<int> main() {
    unusedReturnValue();
}