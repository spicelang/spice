// Std imports
import "std/data/unordered-map";

// Own imports
import "bootstrap/reader/code-loc";
//import "bootstrap/source-file";

type ScopeType enum {
    GLOBAL,
    FUNC_PROC_BODY,
    LAMBDA_BODY,
    STRUCT,
    INTERFACE,
    ENUM,
    IF_ELSE_BODY,
    WHILE_BODY,
    FOR_BODY,
    FOREACH_BODY,
    CASE_BODY,
    DEFAULT_BODY,
    UNSAFE_BODY,
    ANONYMOUS_BLOCK_BODY
}

/**
 * Represents an enclosed group of instructions, which are semantically separated from other scopes.
 * In the source code, scopes usually are written as curly braces.
 *
 * Following language structures use scopes:
 * - global scope
 * - functions/procedures
 * - structs
 * - enums
 * - interfaces
 * - thread blocks
 * - unsafe blocks
 * - for loops
 * - foreach loops
 * - while loops
 * - if statements
 * - anonymous scopes
 */
type Scope struct {
    // Public members
    public Scope* parent
    public SourceFile* sourceFile
    public Map<String, Scope> children
    public SymbolTable symbolTable
    public CodeLoc* codeLoc = nil<CodeLoc*>
    public ScopeType scopeType
    public bool isGenericScope = false
    public bool isAsyncScope = false
    public bool isDtorScope = false
    // Private members
    FunctionRegistry functions
    StructRegistry structs
    InterfaceRegistry interfaces
    UnorderedMap<String, GenericType> genericTypes
}

p Scope.ctor(Scope* parent, SourceFile* sourceFile, ScopeType scopeType, const CodeLoc *codeLoc) {
    this.parent = parent;
    this.sourceFile = sourceFile;
    this.scopeType = scopeType;
    this.symbolTable = SymbolTable(parent == nil<Scope*> ? nil<SymbolTable*> : &parent.symbolTable, this);
    this.codeLoc = codeLoc;
}

/**
 * Create a child scope and return it
 *
 * @param scopeName Name of the child scope
 * @param scopeType Type of the child scope
 * @param declCodeLoc Code location of the scope
 * @return Child scope (heap allocated)
 */
f<Scope*> Scope.createChildScope(const String& scopeName, ScopeType scopeType, const CodeLoc *declCodeLoc) {
    children[scopeName] = Scope(this, sourceFile, scopeType, declCodeLoc);
    return &children[scopeName];
}

/**
 * Rename the child scope. This is useful for realizing function overloading by storing a function with not
 * only its name, but also its signature
 *
 * @param oldName Old name of the child table
 * @param newName New name of the child table
 */
p Scope.renameChildScope(const String& oldName, const String& newName) {
    assert children.contains(oldName) && !children.contains(newName);
    children[newName] = children[oldName];
    children.erase(oldName);
}

/**
 * Duplicates the child scope by copying it. The duplicated symbols point to the original ones.
 *
 * @param oldName Old name of the child block
 * @param newName New block name
 */
p Scope.copyChildScope(const String& oldName, const String& newName) {
    assert children.constains(oldName) && !children.contains(newName);
    // Create copy
    Scope* child = children.at(oldName);
    const heap Scope* newScope = child.deepCopyScope();
    // Save copy under new name
    children[newName] = newScope;
}

/**
 * Deep copy the current scope and all its children
 *
 * @return Deep copy of the current scope
 */
f<heap Scope*> Scope.deepCopyScope() {
    const heap Scope* newScope; // ToDo: Extend
    return newScope;
}

/**
 * Get a child scope of the current scope by its name
 *
 * @param scopeName Child scope name
 * @return Child scope
 */
f<Scope*> Scope.getChildScope(const String& scopeName) {
    if this.children.isEmpty() && this.children.contains(scopeName) {
        return this.children.get(scopeName);
    }
    return nil<Scope*>;
}

/**
 * Retrieve all variables in the current scope, that have reached the end of their lifetime at the end of this scope
 *
 * @return Collection of EOL variables
 */
f<Vector<SymbolTableEntry*>> Scope.getVarsGoingOutOfScope() {
    assert this.parent != nil<Scope*>; // Should not be called in root scope
    Vector<SymbolTableEntry*> varsGoingOutOfScope;

    // Collect all variables in this scope
    foreach const Pair<String, SymbolTableEntry*> symbol : this.symbolTable.symbols {
        const String& name = symbol.getFirst();
        const SymbolTableEntry* entry = symbol.getSecond();
        // Skip 'this' and result variables
        if name == THIS_VARIABLE_NAME || name == RETURN_VARIABLE_NAME {
            continue;
        }
        // Skip parameters (ToDo: Remove when copy constructors work for by-value argument passing)
        if entry.isParam {
            continue;
        }
        // Found variable, that goes out of scope
        varsGoingOutOfScope.push(&this.symbolTable.symbols.get(name));
    }

    // If this is the scope of a dtor, also return all fields of the struct
    if this.isDtorScope {
        assert this.parent != nil<Scope*> && this.parent.scopeType == ScopeType::STRUCT;
        // Get all fields of the struct
        foreach const Pair<String, SymbolTableEntry*> field : paren.symbolTable.symbols {
            const String& name = symbol.getFirst();
            const SymbolTableEntry* entry = symbol.getSecond();
            const QualType& qualType = entry.getQualType();
            if !qualType.isOneOf([TY_FUNCTION, TY_PROCEDURE]) {
                varsGoingOutOfScope.push(&field.getSecond());
            }
        }
    }

    return varsGoingOutOfScope;
}
