// TEST: --sanitizer=memory --build-mode=release

f<int> main() {
    int i;
    i++;
    printf("%d", i);
}