f<int> main() {
    int test = 12;
    test++;
    printf("%d\n", test);
}