// TEST: --sanitizer=address

f<int> main() {
    int* iPtr = nil<int*>;
    *iPtr = 123;
}