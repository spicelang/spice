import "std/runtime/string_rt" as _rt_str;

f<int> main() {
    _rt_str::String s = _rt_str::String("Hello ");
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.append("World!");
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.appendChar('?');
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.appendChar('!');
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    printf("Equals: %d\n", s.opEquals("Hello World!?!"));
    printf("Equals: %d\n", s.opEquals("Hello World!!"));
    printf("Not Equals: %d\n", s.opNotEquals("Hello World!?!"));
    printf("Not Equals: %d\n", s.opNotEquals("Hello World!!"));
    s.clear();
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.reserve(100l);
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d", s.getCapacity());
}