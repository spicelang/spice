/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/data/vector" as vector;

f<int> main() {
    dyn v = vector.Vector<int>{};
    v.push(4);
    v.push(2);
}*/

/*f<int> testFunc(string param = "Test") {
    printf("Test func %s\n", param);
    return 2;
}

f<int> main() {
    int res = testFunc();
    printf("Result: %d\n", res);
}*/

/*type T dyn;
type U dyn;

f<double> genericFunction<T, U>(T arg1, U arg2, int arg3 = 10) {
    return arg1 + arg2 + arg3;
}

f<double> genericFunction<T, U>(T arg1, U arg2, T arg3) {
    return arg1 + arg2 + arg3;
}

f<int> main() {
    printf("%f\n", genericFunction<int, double>(1, 2.4));
    printf("%f\n", genericFunction<long, double>(12l, 2.0));
}*/

import "os-test2" as s1;

f<int> main() {
    //s1.printFormat<double>(1.123);
    //s1.printFormat<int>(543);
    //s1.printFormat<string[]>({"Hello", "World"});
}