import "std/data/linked-list";

f<int> main() {
    LinkedList<int> ll;
    ll.insert(1);
    ll.insert(2);
    ll.insert(3);
    ll.insertAt(3, 1);
}