#[core.linker.dll]
p testFunction() {}

f<int> main() {
    testFunction();
}