import "test-program" as test;