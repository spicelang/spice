// Std imports
import "std/data/vector";

// Own imports
import "bootstrap/model/function-intf";
import "bootstrap/model/struct-intf";
import "bootstrap/model/interface-intf";

// Operator overload function names
public const string OP_FCT_PREFIX = "op.";
public const string OP_FCT_PLUS = "op.plus";
public const string OP_FCT_MINUS = "op.minus";
public const string OP_FCT_MUL = "op.mul";
public const string OP_FCT_DIV = "op.div";
public const string OP_FCT_EQUAL = "op.equal";
public const string OP_FCT_NOT_EQUAL = "op.notequal";
public const string OP_FCT_SHL = "op.shl";
public const string OP_FCT_SHR = "op.shr";
public const string OP_FCT_PLUS_EQUAL = "op.plusequal";
public const string OP_FCT_MINUS_EQUAL = "op.minusequal";
public const string OP_FCT_MUL_EQUAL = "op.mulequal";
public const string OP_FCT_DIV_EQUAL = "op.divequal";
public const string OP_FCT_POSTFIX_PLUS_PLUS = "op.plusplus.post";
public const string OP_FCT_POSTFIX_MINUS_MINUS = "op.minusminus.post";
public const string OP_FCT_SUBSCRIPT = "op.subscript";

/**
 * Saves a constant value for an AST node to realize features like array-out-of-bounds checks
 */
public type CompileTimeValue struct {
    double doubleValue = 0.0
    int intValue = 0
    short shortValue = 0s
    long longValue = 0l
    byte byteValue = (byte) 0
    char charValue = '\0'
    unsigned long stringValueOffset = 0l // Offset into vector of strings in GlobalResourceManager
    bool boolValue = false
}

public type IASTNode interface {
    public f<Vector<IASTNode*>> getChildren();
    public f<Vector<Vector<const IFunction*>>> getOpFctPointers();
    public p customItemsInitialization(unsigned long /*manifestationCount*/);
    public f<bool> hasCompileTimeValue();
    public f<CompileTimeValue> getCompileTimeValue();
    public f<bool> returnsOnAllControlPaths(bool* /*doSetPredecessorsUnreachable*/);
    public f<Vector<IFunction*>*> getFctManifestations(const String&);
    public f<Vector<IStruct*>*> getStructManifestations();
    public f<Vector<IInterface*>*> getInterfaceManifestations();
    public f<bool> isFctOrProcDef();
    public f<bool> isStructDef();
    public f<bool> isParam();
    public f<bool> isStmtLst();
    public f<bool> isAssignExpr();
    public f<bool> isExprStmt();
}