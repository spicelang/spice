//import "std/type/int" as unused;

f<int> main() {
    unsigned int t = 12u;
    printf("%d", t);
}