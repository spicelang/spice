import "std/io/dir" as dir;

f<int> main() {
    dir.listDir(".\\test\\*.*");
}