f<int> main() {
    int i = 12;
    dyn* test = &i;
}