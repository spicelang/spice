int TEST1 = 10;
string TEST2 = "test string";
double TEST3 = 5.83;
bool TEST4 = false;

f<int> main() {
    TEST1 = 11;
    TEST2 = "test";
    TEST3 = 5.84;
    TEST4 = true;
    printf("Variable values: %d, %s, %f, %u", TEST1, TEST2, TEST3, TEST4);
}