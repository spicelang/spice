public f<String> getLastFragment(String &haystack, const string needle) {
    const unsigned long index = haystack.rfind(needle);
    if index == -1l {
        return haystack;
    }
    return haystack.getSubstring(index + getRawLength(needle));
}