/*import "std/text/print" as print;

type Test struct {
    int field1
    double field2
}

p Test.setField1(int value) {
    this.field1 = value;
}

f<int> Test.getField1() {
    return this.field1;
}

f<int> main() {
    Test test = new Test { 5, 4.567 };
    test.setField1(6);
    print.println("Output:");
    printf("%d", test.getField1());
}*/

f<int> fib(int n) {
    if n <= 2 { return 1; }
    return fib(n - 1) + fib(n - 2);
}

f<int> main() {
    printf("Result: %d", fib(46));
}