import "std/os/os";

import "SourceFile";
import "CliInterface";
import "global/GlobalResourceManager";

/**
 * Compile main source file. All files, that are included by the main source file will be resolved recursively.
 *
 * @param cliOptions Command line options
 * @return Successful or not
 */
f<bool> compileProject(const CliOptions& cliOptions) {
    // Instantiate GlobalResourceManager
    dyn resourceManager = GlobalResourceManager(options);

    // Create source file instance for main source file
    SourceFile* mainSourceFile = resourceManager.createSourceFile(nullptr, MAIN_FILE_NAME, cliOptions.mainFile, false);

    // Run compile pipeline for main source file. All dependent source files are triggered by their parents
    mainSourceFile.runFrontEnd();
    mainSourceFile.runMiddleEnd();
    mainSourceFile.runBackEnd();

    // Link the target executable (link object files to executable)
    resourceManager.linker.prepare();
    resourceManager.linker.link();

    // Print compiler warnings
    mainSourceFile.collectAndPrintWarnings();

    // Print compiler warnings
    mainSourceFile.collectAndPrintWarnings();

    return true;
}

/**
 * Entry point to the Spice compiler
 *
 * @param argc Argument count
 * @param argv Argument vector
 * @return Return code
 */
f<int> main(int argc, string[] argv) {
    // Initialize command line parser
    CliInterface cli;
    cli.create();
    const int exitCode = cli.parse(argc, argv);
    if exitCode != EXIT_SUCCESS {
        return exitCode;
    }

    // Cancel here if we do not have to compile
    if !cli.shouldCompile {
        return EXIT_SUCCESS;
    }

    cli.enrich(); // Prepare the cli options

    // Kick off the compiling process
    if !compileProject(cli.cliOptions) {
        return EXIT_FAILURE;
    }

    // Execute
    if cli.cliOptions.execute {
        cli.runBinary();
    }

    return EXIT_SUCCESS;
}