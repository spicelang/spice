// Imports

public type Generator struct {

}