f<int> main() {
    int i = 123;
    unsigned long j = cast<unsigned long>(i);
    j++;
    printf("i, j: %d, %d", i, j);
}