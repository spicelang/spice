public const unsigned int BYTE_SIZE = 8;
public const unsigned int BYTE_MIN_VALUE = 0;
public const unsigned int BYTE_MAX_VALUE = 255;

// External functions
ext f<unsigned int> snprintf(char*, unsigned long, string, byte);

// Converts a byte to a double
public f<double> toDouble(byte input) {
    return 0.0 + ((int) input);
}

// Converts a byte to an int
public f<int> toInt(byte input) {
    return (int) input;
}

// Converts a byte to a short
public f<short> toShort(byte input) {
    return (short) ((int) input);
}

// Converts a byte to a long
public f<long> toLong(byte input) {
    return (long) ((int) input);
}

// Converts a byte to a char
public f<char> toChar(byte input) {
    return (char) input;
}

// Converts a byte to a string
public f<String> toString(byte input) {
    const unsigned int length = snprintf(nil<char*>, 0l, "%hhu", input);
    result = String(length);
    snprintf((char*) result.getRaw(), length + 1l, "%hhu", input);
}

// Converts a byte to a bool
public f<bool> toBool(byte input) {
    return input == (byte) 1;
}