f<int> main() {
    while true {
        continue 0;
    }
}