f<int> main() {
    p(int, int) add = (int x, int y) -> {
        return x + y;
    };
}