import "std/os/file" as file;

f<int> main() {
    //file.createFile("demo.txt");
    dyn fp = file.openFile("demo.txt", file.MODE_READ_WRITE);
    //printf("FP: %p\n", fp.ptr);
    int r1 = fp.writeChar(65);
    printf("R1: %d\n", r1);
    int r2 = fp.closeFile();
    printf("R2: %d\n", r2);
}