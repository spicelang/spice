import "std/data/set";

f<int> main() {
    Set<int> set;

    // Iterate over empty container
    {
        foreach const int& item : set {
            printf("%d\n", item);
        }
    }

    set.insert(1);
    set.insert(2);
    set.insert(3);
    set.insert(4);
    set.insert(5);
    set.insert(99);
    set.insert(100);
    set.insert(1265);
    set.insert(101);
    set.insert(102);

    // Iterate over filled container
    foreach const int& item : set {
        printf("%d\n", item);
    }
}