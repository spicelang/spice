import "std/data/hash-table";
import "std/data/pair";

f<int> main() {
    HashTable<int, int> table;

    // Iterate over empty container
    {
        foreach Pair<int&, int&> item : table {
            printf("%d: %d\n", item.getFirst(), item.getSecond());
        }
    }

    table.upsert(1, 2);
    table.upsert(2, 3);
    table.upsert(3, 4);
    table.upsert(4, 5);
    table.upsert(5, 6);
    table.upsert(99, 99);
    table.upsert(100, 100);
    table.upsert(1265, 100);
    table.upsert(101, 101);
    table.upsert(102, 102);

    // Iterate over filled container
    foreach Pair<int&, int&> item : table {
        printf("%d: %d\n", item.getFirst(), item.getSecond());
    }
}