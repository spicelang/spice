type TestStruct struct {
    long f1
    int f2
    TestStruct* f3
}

f<int> main() {
    TestStruct ts;
}

/*type TestStruct struct {
    int a = 123
    short b = 1s
}

f<int> main() {
    TestStruct ts;
    printf("%d %d\n", ts.a, ts.b);
}*/