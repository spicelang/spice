/**
 * Check if an int is a power of two
 *
 * @param input Input number
 * @return Is power of two
 */
public f<bool> isPowerOfTwo(int input) {
    return (input & (input - 1)) == 0;
}