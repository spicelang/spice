import "std/io/cli-parser";

type CliOptions struct {
    bool sayHi = false
}

p callback(bool& value) {
    printf("Callback called with value %d\n", value);
}

f<int> main(int argc, string[] argv) {
    CliParser parser = CliParser("Test Program", "This is a simple test program");
    parser.setVersion("v0.1.0");
    parser.setFooter("Copyright (c) Marc Auberer 2021-2023");

    CliOptions options;
    parser.addFlag("--hi", options.sayHi, "Say hi to the user");
    parser.addFlag("--callback", callback, "Call a callback function");
    parser.addFlag("-cb", p(bool& value) {
        printf("CB called with value %d\n", value);
    }, "Call a callback function");

    parser.parse(argc, argv);

    // Print hi if requested
    if options.sayHi {
        printf("Hi!\n");
    }
}

/*import "std/data/stack";

f<int> main() {
    Stack<int> s1 = Stack<int>{};
    s1.ctor();
    s1.push(123);
    s1.push(456);
    s1.push(789);
    printf("Stack size: %d\n", s1.getSize());
    printf("Stack capacity: %d\n", s1.getCapacity());
    printf("Stack item 3: %d\n", s1.pop());
    printf("Stack item 2: %d\n", s1.pop());
    printf("Stack item 1: %d\n", s1.pop());
}*/

/*type TestStruct struct {
    int a = 123
    short b = 1s
}

f<int> main() {
    TestStruct ts;
    printf("%d %d\n", ts.a, ts.b);
}*/