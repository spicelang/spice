type Stamp struct {
    double value
    bool glued
}

p Stamp.print() {
    printf("Value: %f, glued: %d", this.value, this.glued);
}

type Letter struct {
    string content
    Stamp stamp
}

f<string> Letter.getContent() {
    return this.content;
}

p Letter.setContent(string text) {
    this.content = text;
}

f<Stamp> Letter.getStamp() {
    return this.stamp;
}

p Letter.setStamp(Stamp stamp) {
    this.stamp = stamp;
}

f<int> main() {
    dyn letter = Letter{ "", Stamp{ 3.4, false } };
    printf("Stamp glued: %f\n", letter.getStamp().value);
    letter.getStamp().print();
}

/*import "std/runtime/string_rt" as _rt_str;

f<int> main() {
    printf("%d", _rt_str::String("Test").isEmpty());
}*/

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

/*public f<bool> src(bool x, bool y) {
    return ((x ? 1 : 4) & (y ? 1 : 4)) == 0;
}

public f<int> tgt(int x, int y) {
    return x ^ y;
}

f<int> main() {
    printf("Result: %d, %d", src(false, true), tgt(0, 1));
}*/