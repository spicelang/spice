// Link external functions
ext f<int> getpid();
ext f<int> system(string);

/**
 * Retrieve the process id of the current process.
 *
 * @return Process id
 */
public f<int> getPID() {
    return getpid();
}

/**
 * Executes a shell command by creating a new process.
 *
 * @return Return code of the shell comand
 */
public f<int> execCmd(string cmd) {
    return system(cmd);
}