ext<string> getenv(string);
ext<int> putenv(string);

/**
 * Returns the content of an environment variable as string.
 *
 * @return Env variable content
 */
public f<string> getEnv(string name) {
    return getenv(name);
}

/**
 * Sets the content of an environment variable to the given value.
 *
 * @return Result code: 0 = successful, -1 = failed
 */
public f<int> setEnv(string name, string value) {
    String str = String(name);
    str += "=";
    str += value;
    return putenv(str.getRaw());
}