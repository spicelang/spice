import "source1";

f<int> main() {
    Size test = 23l;
}