/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*f<int> makePi() {
    // Initialize variables
    int q = 1;
    int r = 0;
    int t = 1;
    int k = 1;
    int m = 3;
    int x = 3;
    // Loop
    //int[1000] output = {};
    int outputCounter = 0;
    for int i = 0; i < 1000; i++ {
        if (4 * q + r - t < m * t) {
            //output[outputCounter] = m;
            outputCounter++;
            q = 10 * q;
            r = 10 * (r - m * t);
            t = t;
            k = k;
            m = (10 * (3 * q + r)) / t - 10 * m;
            x = x;
        } else {
            q = q * k;
            r = (2 * q + r) * x;
            t = t * x;
            k = k + 1;
            m = (q * (7 * k + 2) + r * x) / (t * x);
            x = x + 2;
        }
    }
    return 3;
}

f<int> main() {
    makePi();
}*/

/*import "std/io/dir" as dir;

f<int> main() {
    dir.mkDir("./test", dir.MODE_ALL_RWX);
}*/





/*const int AF_INET = 2;
const int SOCK_STREAM = 1;
const int IPPROTO_IP = 0;

type InAddr struct {
    unsigned int addr
}

type SockAddrIn struct {
    unsigned short sinFamily
    unsigned short sinPort
    InAddr sinAddr
}

type Socket struct {
    int sockFd // Actual socket
    int connFd // Current connection
    short errorCode
}

ext<int> socket(int, int, int);
ext<int> accept(int, SockAddrIn*, int);

f<int> Socket.acceptConnection() {
    SockAddrIn cliAddr = SockAddrIn {};
    this.connFd = accept(this.sockFd, &cliAddr, 16);
    if this.connFd == -1 {
        //result.errorCode = ERROR_ACCEPT;
        return -1;
    }
    return this.connFd;
}

f<int> openServerSocket(unsigned short port) {
    Socket s = Socket { socket(AF_INET, SOCK_STREAM, IPPROTO_IP), 0, 0s };

    s.acceptConnection();

    return s.sockFd;
}

f<int> main() {
    openServerSocket(8080s);
}*/




const int AF_INET = 2;
const int SOCK_STREAM = 1;
const int SOCK_DGRAM = 2;
const int IPPROTO_IP = 0;
const int IPPROTO_UDP = 17;
const int INADDR_ANY = 0;

type InAddr struct {
    unsigned int addr
}

type SockAddrIn struct {
    unsigned short sinFamily
    unsigned short sinPort
    InAddr sinAddr
}

type Socket struct {
    int sockFd // Actual socket
    int connFd // Current connection
    short errorCode
}

const short ERROR_SOCKET = -1s;
const short ERROR_BIND = -2s;
const short ERROR_LISTEN = -3s;
const short ERROR_ACCEPT = -4s;

ext<int> socket(int, int, int);
ext<int> bind(int, SockAddrIn*, int);
ext<int> listen(int, int);
ext<int> accept(int, SockAddrIn*, int);
ext<int> close(int);
ext<int> htonl(int);     // Fairly simple to re-implement in Spice
ext<short> htons(short); // Fairly simple to re-implement in Spice

/**
 * Accept an incoming connection to the socket and save the connection file desceiptor
 * to the socket object.
 *
 * @return Connection file descriptor
 */
f<int> Socket.acceptConnection() {
    SockAddrIn cliAddr = SockAddrIn {};
    this.connFd = accept(this.sockFd, &cliAddr, 16 /* hardcoded sizeof(cliAddr) */);
    if this.connFd == -1 {
        //result.errorCode = ERROR_ACCEPT;
        return -1;
    }
    return this.connFd;
}

p Socket.waitForIncomingConnections() {
    // ToDo: Implement
}

/**
 * Closes the socket. This method should always be called by the user before exiting the program.
 *
 * @return Error code for closing the socket
 */
f<int> Socket.close() {
    return close(this.sockFd);
}

f<int> openServerSocket(unsigned short port) {
    Socket s = Socket { socket(AF_INET, SOCK_STREAM, IPPROTO_IP), 0, 0s };

    // Cancel on failure
    if s.sockFd == -1 {
        //result.errorCode = ERROR_SOCKET;
        return -1;
    }

    InAddr inAddr = InAddr { htonl(INADDR_ANY) };
    SockAddrIn servaddr = SockAddrIn { (short) AF_INET, htons(port), inAddr };

    int bindResult = bind(s.sockFd, &servaddr, 16 /* hardcoded sizeof(servaddr) */);
    if bindResult != 0 {
        //result.errorCode = ERROR_BIND;
        return -2;
    }

    int listenResult = listen(s.sockFd, 5 /* backlog */);
    if listenResult != 0 {
        //result.errorCode = ERROR_LISTEN;
        return -3;
    }

    s.acceptConnection();

    return s.sockFd;
}

// Tmp function until bug #95 is fixed
f<int> closeSocket(int fd) {
    return close(fd);
}

f<int> main() {
    openServerSocket(8080s);
}