import "std/runtime/string" as str;

f<int> main() {
    string a = "Hello ";
    string b = "World!";
    printf("String a: %s", a);
    printf("String b: %s", b);
    //printf("String a+b: %s", a + b);
}