public const int SIZE = 64;
public const long MIN_VALUE = -9223372036854775808l;
public const long MAX_VALUE = 9223372036854775807l;

const int nSmall = 100;
const string smallsString10 = "0123456789";
const string smallsString100 = "00010203040506070809101112131415161718192021222324252627282930313233343536373839404142434445464748495051525354555657585960616263646566676869707172737475767778798081828384858687888990919293949596979899";

// Converts a long to a double
public f<double> toDouble(long input) {
    return 0.0 + input;
}

// Converts a long to an int
public f<int> toInt(long input) {
    return (int) input;
}

// Converts a long to a short
public f<short> toShort(long input) {
    return (short) input;
}

// Converts a long to a byte
public f<byte> toByte(long input) {
    return (byte) ((int) input);
}

// Converts a long to a char
public f<char> toChar(long input) {
    return (char) input;
}

// Converts a long to a string
public f<string> toString(long input) {
    // ToDo: Implement (See https://github.com/golang/go/blob/master/src/strconv/itoa.go)
    return "";
}

// Converts a long to a boolean
public f<bool> toBool(long input) {
    return input >= 1;
}

// Check if the input is a power of two
public f<bool> isPowerOfTwo(long input) {
    return (input & (input - 1l)) == 0l;
}