// Std imports
import "std/data/vector";
import "std/data/map";

// Helper structs
public type Param struct {
    Type sType
    bool isOptional
}

public type NamedParam struct {
    String name
    Type sType
    bool isOptional
}

// Type aliases
type ParamList alias Vector<Param>;
type NamedParamList alias Vector<NamedParam>;

public type Function struct {
    String name
    Type thisType
    Type returnType
    ParamLits paramList
    Vector<GenericType> templateTypes
    Map<String, Type> typeMapping
    SymbolTableEntry* entry
    ASTNode* declNode
    bool genericSubstantiation
    bool alreadyTypeChecked
    bool external
    bool used
}