type T dyn;

f<int> main() {
    printf("Alignment: %d", alignof(T));
}