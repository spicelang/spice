import "std/iterator/iterable";
import "std/data/pair";

type MockIterator struct : Iterable<int> {
    int item
    unsigned long cursor
}

p MockIterator.ctor() {
    this.cursor = 0l;
}

f<int&> MockIterator.get() {
    return this.item;
}

f<Pair<unsigned long, int&>> MockIterator.getIdx() {
    return Pair<unsigned long, int&>(0l, this.item);
}

f<bool> MockIterator.isValid() {
    return true;
}

p MockIterator.next() {}

f<int> main() {
    foreach dyn demoItem : MockIterator() {
        printf("Demo item\n");
    }
}