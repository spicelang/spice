import "std/data/hash-table";

f<int> main() {
    HashTable<int, int> hashTable = HashTable<int, int>();
    hashTable.upsert(1, 2);
    hashTable.upsert(2, 3);

    Optional<int> value = hashTable.get(1);
    assert(value.get() == 2);
    value = hashTable.get(2);
    assert(value.get() == 3);

}

/*import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

f<int> main() {
    DefaultMemoryManager defaultMemoryManager;
    IMemoryManager* memoryManager = &defaultMemoryManager;
    BlockAllocator<int> allocator = BlockAllocator<int>(memoryManager, 10l);
}*/