f<string> getOsName() {
    return "windows";
}