import "std/data/vector";

f<int> main() {
    Vector<String> vec;
    vec.pushBack(String("Hello"));
    vec.pushBack(String("Dear"));
    vec.pushBack(String("\n World"));

    vec[1][2] = 'p';
    String& item0 = vec[0];
    item0.replaceAll("l", "x");
    String& item2 = vec.get(2);
    item2 = item2.trim();

    foreach String s : vec {
        printf("%s\n", s);
    }
}