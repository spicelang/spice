import "std/data/vector";

f<Vector<string>> getStringVec() {
    Vector<string> queue;
    queue.pushBack("Hello");
    queue.pushBack("World");
    return queue;
}

f<int> main() {
    const Vector<string> args = getStringVec();
    foreach unsigned long i, const string& arg : args {
        printf("Arg %d: %s\n", i, arg);
    }
}