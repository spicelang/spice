f<int> main() {
    if (1 == 1) {
        printf("Test: %s", "Value");
    }
    return 0;
}