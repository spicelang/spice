// See Issue #155 (fixed)

type T dyn;

public type Vector<T> struct {
    T* contents
    unsigned long capacity
    unsigned long size
    unsigned int itemSize
}

public f<int> Vector.get(long index) {
    if (index <= size) { // size instead this.size
        return 1;
    }
    return 0;
}

f<int> main() {
    dyn v = Vector<int>{};
    int v0 = v.get(0l);
}