type TestStruct struct {
    int field
}

f<int> main() {
    printf("Size: %d", sizeof(TestStruct));
}