import "std/io/csv";
import "std/io/filepath";

type Row struct : CSVRow {
    string name
    int age
    string city
    double salary
}

f<int> main() {
    FilePath filePath = FilePath("/home/marc/Documents/Dev/spice/test/test-files/std/io/csv-parser/input.csv");
    CSVParser<Row> parser = CSVParser<Row>(filePath, ',');
    CSVTable<Row> table = parser.parse();
    // Print the headers
    printf("Headers: ");
    for unsigned long i = 0l; i < table.headers.getSize(); i++ {
        printf("%s, ", table.headers[i]);
    }
}
