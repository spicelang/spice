import "std/type/type-conversion";
import "std/type/short";

f<int> main() {
    // toDouble()
    double asDouble = toDouble(123s);
    assert asDouble == 123.0;

    // toInt()
    int asInt = toInt(-345s);
    assert asInt == -345;

    // toLong()
    long asLong = toLong(45s);
    assert asLong == 45l;

    // toByte()
    byte asByte = toByte(12s);
    assert asByte == cast<byte>(12);

    // toChar()
    char asChar = toChar(66s);
    assert asChar == 'B';

    // toString()
    String asString = toString(15s);
    assert asString.getRaw() == "15";

    // toBool()
    bool asBool1 = toBool(1s);
    assert asBool1 == true;
    bool asBool2 = toBool(0s);
    assert asBool2 == false;

    // isPowerOfTwo()
    assert isPowerOfTwo(16s);
    assert !isPowerOfTwo(31s);

    printf("All assertions succeeded");
}