// Imports
import "std/text/print";
import "std/data/pair";
import "CliInterface";
import "ast/AstNodes";

type CompileStageType enum {
    NONE,
    LEXER,
    PARSER,
    CST_VISUALIZER,
    AST_BUILDER,
    AST_OPTIMIZER,
    AST_VISUALIZER,
    IMPORT_COLLECTOR,
    SYMBOL_TABLE_BUILDER,
    TYPE_CHECKER_PRE,
    TYPE_CHECKER_POST,
    BORROW_CHECKER,
    ESCAPE_ANALYZER,
    IR_GENERATOR,
    IR_OPTIMIZER,
    OBJECT_EMITTER
}

type CompileStageIOType enum {
    IO_CODE,
    IO_TOKENS,
    IO_CST,
    IO_AST,
    IO_IR,
    IO_OBJECT_FILE
}

type TimerOutput struct {
  unsigned long lexer = 0
  unsigned long parser = 0
  unsigned long cstVisualizer = 0
  unsigned long astBuilder = 0
  unsigned long astOptimizer = 0
  unsigned long astVisualizer = 0
  unsigned long importCollector = 0
  unsigned long symbolTableBuilder = 0
  unsigned long typeCheckerPre = 0
  unsigned long typeCheckerPost = 0
  unsigned long borrowChecker = 0
  unsigned long escapeAnalyzer = 0
  unsigned long irGenerator = 0
  unsigned long irOptimizer = 0
  unsigned long objectEmitter = 0
  unsigned long executionEngine = 0
}

/**
 * Collects the output of the compiler for debugging
 */
type CompilerOutput struct {
    String cstString
    String astString
    String symbolTableString
    String irString
    String irOptString
    String asmString
    Vector<CompilerWarning> warnings
    TimerOutput times
}

type NameRegistryEntry struct {
    String name
    SymbolTableEntry* targetEntry
    Scope* targetScope
    SymbolTableEntry* importEntry
    String predecessorName
}

/**
 * Represents a single source file
 */
public type SourceFile struct {
    public String name
    public String fileName
    public String filePath
    public String fileDir
    public String objectFilePath
    public bool stdFile = false
    public bool mainFile = true
    public CompilerOutput compilerOutput
    public SourceFile* parent
    public String cacheKey
    public bool restoredFromCache = false
    public EntryNode ast
    public Scope globalScope
    //public llvm::Module llvmModule
    public Map<String, Pair<SourceFile, const ASTNode*>> dependencies
    public Map<String, NameRegistryEntry> exportedNameRegistry

    GlobalResourceManager& resourceManager
    unsigned short importedRuntimeModules = 0
    unsigned short typeCheckerRuns = 0
}

public p SourceFile.ctor(GlobalResourceManager &resourceManager, SourceFile* parent, string name, string filePath, bool stdFile) {
    // Copy data
    this.resourceManager = resourceManager;
    this.parent = parent;
    this.name = name;
    this.filePath = filePath;
    this.stdFile = stdFile;

    // Deduce fileName and fileDir
    /*this.fileName = ;
    this.fileDir = ;*/
}

public p SourceFile.runLexer() {
    // Lex this source file
}

public p SourceFile.runParser() {
    // Parse this source file
}

public p SourceFile.runCSTVisualizer(string* output) {
    // Only execute if enabled
    if !cliOptions.dumpCST && !cliOptions.testMode { return; }

    // ToDo: Extend
}

public p SourceFile.runASTBuilder() {
    // Transform the imported source files
    // ToDo: Extend
}

public p SourceFile.runASTVisualizer(string* output) {
    // Only execute if enabled
    if !cliOptions.dumpAST && !cliOptions.testMode { return; }

    // ToDo: Extend
}

public p SourceFile.runImportCollector() {

}

public p SourceFile.runSymbolTableBuilder() {

}

public p SourceFile.runTypeChecker() {

}

p SourceFile.runTypeCheckerPre() {

}

p SourceFile.runTypeCheckerPost() {

}

public p SourceFile.runBorrowChecker() {

}

public p SourceFile.runEscapeAnalyzer() {

}

public p SourceFile.runIRGenerator() {

}

public p SourceFile.runDefaultIROptimizer() {

}

public p SourceFile.runObjectEmitter() {

}

public p SourceFile.concludeCompilation() {

}

public f<int> SourceFile.execute() {

}

public p SourceFile.runFrontEnd() {

}

public p SourceFile.runMiddleEnd() {

}

public p SourceFile.runBackEnd() {

}

f<bool> SourceFile.isAlreadyImported(const string filePathSearch) {
    // Check if the current source file corresponds to the path to search
    if filePath == filePathSearch { return true; }
    // Check parent recursively
    return parent != nil<SourceFile*> && parent.isAlreadyImported(filePathSearch);
}