type T int|long|short;

type Compareable<T> interface {
    f<T**> compare();
}

f<int> main() {

}