unsigned short UNSIGNED_SHORT = -10;
const signed int TEST = 6s;

f<int> main() {
    printf("Int: %d", TEST);
}