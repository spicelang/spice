f<int> main() {
    Test inst = new Test { false };
    printf("%u", inst.testField);
}

type Test struct {
    bool testField
}