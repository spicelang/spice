f<int> main() {
    short**[8] _ = {};
}