f<int> main() {
    int& ref;
}