// Link WinSock library
#![core.linux.linker.flag = "-lws2_32"]

// Import common logic
import "std/net/socket";

const unsigned short REQUESTED_WSA_VERSION = 514s;

type WSAData struct {
    unsigned short wVersion
    unsigned short wHighVersion
    unsigned short iMaxSockets
    unsigned short iMaxUdpDg
    char* lpVendorInfo
    char[257] szDescription
    char[129] szSystemStatus
}

ext f<int> WSAStartup(short, WSAData*);
ext f<int> WSACleanup();
ext f<int> socket(int, int, int);
ext f<int> bind(int, SockAddrIn*, unsigned int);
ext f<int> listen(int, int);
ext f<int> accept(int, SockAddrIn*, unsigned int);
ext f<int> close(int);
ext f<int> htonl(int);     // Fairly simple to re-implement in Spice
ext f<short> htons(short); // Fairly simple to re-implement in Spice

public type Socket struct {
    int sockFd // Actual socket
    int connFd // Current connection
}

public p Socket.dtor() {
    this.close();
}

/**
 * Accept an incoming connection to the socket and save the connection file desceiptor
 * to the socket object.
 *
 * @return Connection file descriptor
 */
public f<Result<int>> Socket.acceptConnection() {
    SockAddrIn cliAddr = SockAddrIn {};
    this.connFd = accept(this.sockFd, &cliAddr, (unsigned int) sizeof(cliAddr));
    if this.connFd == -1 {
        return err<int>(Error("Error while accepting connection"));
    }
    return ok(this.connFd);
}

/**
 * Closes the socket. This method should always be called by the user before exiting the program.
 *
 * @return Closing the connection was successful or not
 */
public f<bool> Socket.close() {
    return close(this.sockFd) == 0 && WSACleanup() == 0;
}

/**
 * Opens a TCP server socket and exposes it to the given port.
 * The maxWaitingConnections defines the maximum length to which the queue of pending connections may grow. If a
 * connection request arrives when the queue is full, the client may receive an error with an indication of
 * ECONNREFUSED or, if the underlying protocol support retransmission, the request may be ignored so that a later
 * reattempt at connection succeeds.
 *
 * @param port Port to open the socket on
 * @param maxWaitingConnections Maximum size of the queue of pending client connections
 * @return Socket file descriptor
 */
public f<Result<Socket>> openServerSocket(unsigned short port, int maxWaitingConnections = 5) {
    WSAData wsaData = WSAData{};
    if WSAStartup(REQUESTED_WSA_VERSION, &wsaData) != 0 {
        return err<Socket>(Error("Error initializing WSA"));
    }

    const Socket s = Socket { socket(AF_INET, SOCK_STREAM, IPPROTO_IP), 0 };

    // Cancel on failure
    if s.sockFd == -1l {
        return err<Socket>(Error("Error creating socket"));
    }

    InAddr inAddr = InAddr { htonl(INADDR_ANY) };
    SockAddrIn servAddr = SockAddrIn { (short) AF_INET, htons(port), inAddr };

    int bindResult = bind(s.sockFd, &servAddr, (unsigned int) sizeof(servAddr));
    if bindResult != 0 {
        return err<Socket>(Error("Error binding to address"));
    }

    int listenResult = listen(s.sockFd, maxWaitingConnections);
    if listenResult != 0 {
        return err<Socket>(Error("Error listening on address"));
    }

    s.acceptConnection();

    return ok(s);
}
