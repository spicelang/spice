type TLhs dyn;
type TRhs dyn;
type TRes dyn;

// ------------------------------------------ += ------------------------------------------

p plusEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs += rhs;
    assert lhs == expectedResult;
}

p plusEqualTestInnerUnsafe<TRhs>(int* lhs, const TRhs rhs, const int* expectedResult) {
    unsafe {
        lhs += rhs;
    }
    assert lhs == expectedResult;
}

p plusEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    plusEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    plusEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    plusEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    plusEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p plusEqualTest() {
    // Lhs is double
    plusEqualTestOuter<double, double>(1.234, 98.7654, 99.9994, -99.9994, 97.5314, -97.5314);
    // Lhs is int
    plusEqualTestOuter<int, int>(78, 674, 752, -752, 596, -596);
    plusEqualTestOuter<int, short>(78, 7s, 85, -85, -71, 71);
    plusEqualTestOuter<int, long>(78, 2384723l, 2384801, -2384801, 2384645, -2384645);
    // Lhs is short
    plusEqualTestOuter<short, int>(78s, 674, 752s, -752s, 596s, -596s);
    plusEqualTestOuter<short, short>(78s, 7s, 85s, -85s, -71s, 71s);
    plusEqualTestOuter<short, long>(78s, 2384723l, 25505s, -25505s, 25349s, -25349s);
    // Lhs is long
    plusEqualTestOuter<long, int>(78l, 674, 752l, -752l, 596l, -596l);
    plusEqualTestOuter<long, short>(78l, 7s, 85l, -85l, -71l, 71l);
    plusEqualTestOuter<long, long>(78l, 2384723l, 2384801l, -2384801l, 2384645l, -2384645l);
    // Lhs is char
    plusEqualTestInner<char, int>('A', 5, 'F');
    plusEqualTestInner<char, int>('A', -5, '<');
    // Lhs is ptr
    int[5] input = [0, 0, 0, 0, 0];
    plusEqualTestInnerUnsafe(&input[2], 2, &input[4]);
    plusEqualTestInnerUnsafe(&input[2], -2, &input[0]);
    plusEqualTestInnerUnsafe(&input[2], 2s, &input[4]);
    plusEqualTestInnerUnsafe(&input[2], -2s, &input[0]);
    plusEqualTestInnerUnsafe(&input[2], 2l, &input[4]);
    plusEqualTestInnerUnsafe(&input[2], -2l, &input[0]);
}

// ------------------------------------------ -= ------------------------------------------

p minusEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs -= rhs;
    assert lhs == expectedResult;
}

p minusEqualTestInnerUnsafe<TRhs>(int* lhs, const TRhs rhs, const int* expectedResult) {
    unsafe {
        lhs -= rhs;
    }
    assert lhs == expectedResult;
}

p minusEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    minusEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    minusEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    minusEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    minusEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p minusEqualTest() {
    // Lhs is double
    minusEqualTestOuter<double, double>(1.234, 98.7654, -97.5314, 97.5314, -99.9994, 99.9994);
    // Lhs is int
    minusEqualTestOuter<int, int>(78, 674, -596, 596, -752, 752);
    minusEqualTestOuter<int, short>(78, 7s, 71, -71, -85, 85);
    minusEqualTestOuter<int, long>(78, 2384723l, -2384645, 2384645, -2384801, 2384801);
    // Lhs is short
    minusEqualTestOuter<short, int>(78s, 674, -596s, 596s, -752s, 752s);
    minusEqualTestOuter<short, short>(78s, 7s, 71s, -71s, -85s, 85s);
    // Note: wrap-around consistent with short semantics
    minusEqualTestOuter<short, long>(78s, 2384723l, cast<short>(78s - 2384723l), cast<short>(-78s - -2384723l), cast<short>(-78s - 2384723l), cast<short>(78s - -2384723l));
    // Lhs is long
    minusEqualTestOuter<long, int>(78l, 674, -596l, 596l, -752l, 752l);
    minusEqualTestOuter<long, short>(78l, 7s, 71l, -71l, -85l, 85l);
    minusEqualTestOuter<long, long>(78l, 2384723l, -2384645l, 2384645l, -2384801l, 2384801l);
    // Lhs is char
    minusEqualTestInner<char, int>('A', 5, '<');
    minusEqualTestInner<char, int>('A', -5, 'F');
    // Lhs is ptr
    int[5] input = [0, 0, 0, 0, 0];
    minusEqualTestInnerUnsafe(&input[2], 2, &input[0]);
    minusEqualTestInnerUnsafe(&input[2], -2, &input[4]);
    minusEqualTestInnerUnsafe(&input[2], 2s, &input[0]);
    minusEqualTestInnerUnsafe(&input[2], -2s, &input[4]);
    minusEqualTestInnerUnsafe(&input[2], 2l, &input[0]);
    minusEqualTestInnerUnsafe(&input[2], -2l, &input[4]);
}

// ------------------------------------------ *= ------------------------------------------

p mulEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs *= rhs;
    assert lhs == expectedResult;
}

p mulEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    mulEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    mulEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    mulEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    mulEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p mulEqualTest() {
    // Lhs double
    mulEqualTestOuter<double, double>(1.5, 2.0, 3.0, 3.0, -3.0, -3.0);
    // Lhs int
    mulEqualTestOuter<int, int>(6, 7, 42, 42, -42, -42);
    mulEqualTestOuter<int, short>(6, 3s, 18, 18, -18, -18);
    mulEqualTestOuter<int, long>(6, 5l, 30, 30, -30, -30);
    // Lhs short
    mulEqualTestOuter<short, int>(6s, 7, 42s, 42s, -42s, -42s);
    mulEqualTestOuter<short, short>(6s, 3s, 18s, 18s, -18s, -18s);
    // Note: wrap-around consistent with short semantics
    mulEqualTestOuter<short, long>(200s, 2000l, cast<short>(200 * 2000), cast<short>(-200 * -2000), cast<short>(-200 * 2000), cast<short>(200 * -2000));
    // Lhs long
    mulEqualTestOuter<long, int>(6l, 7, 42l, 42l, -42l, -42l);
    mulEqualTestOuter<long, short>(6l, 3s, 18l, 18l, -18l, -18l);
    mulEqualTestOuter<long, long>(6l, 5l, 30l, 30l, -30l, -30l);
}

// ------------------------------------------ /= ------------------------------------------

p divEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs /= rhs;
    assert lhs == expectedResult;
}

p divEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    divEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    divEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    divEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    divEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p divEqualTest() {
    // Lhs double
    divEqualTestOuter<double, double>(9.0, 3.0, 3.0, 3.0, -3.0, -3.0);
    // Lhs int
    divEqualTestOuter<int, int>(42, 7, 6, 6, -6, -6);
    divEqualTestOuter<int, short>(42, 3s, 14, 14, -14, -14);
    divEqualTestOuter<int, long>(42, 6l, 7, 7, -7, -7);
    // Lhs short
    divEqualTestOuter<short, int>(42s, 7, 6s, 6s, -6s, -6s);
    divEqualTestOuter<short, short>(42s, 3s, 14s, 14s, -14s, -14s);
    divEqualTestOuter<short, long>(100s, 25l, 4s, 4s, -4s,- 4s);
    // Lhs long
    divEqualTestOuter<long, int>(42l, 7, 6l, 6l, -6l, -6l);
    divEqualTestOuter<long, short>(42l, 3s, 14l, 14l, -14l, -14l);
    divEqualTestOuter<long, long>(42l, 6l, 7l, 7l, -7l, -7l);
}

// ------------------------------------------ %= ------------------------------------------

p remEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs %= rhs;
    assert lhs == expectedResult;
}

p remEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    remEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    remEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    remEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    remEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p remEqualTest() {
    // Lhs double
    remEqualTestOuter<double, double>(9.0, 3.0, 0.0, 0.0, 0.0, 0.0);
    // Lhs int
    remEqualTestOuter<int, int>(42, 7, -0, -0, 0, 0);
    remEqualTestOuter<int, short>(42, 8s, 2, -2, -2, 2);
    remEqualTestOuter<int, long>(42, 9l, 6, -6, -6, 6);
    // Lhs short
    remEqualTestOuter<short, int>(42s, 7, -0s, -0s, 0s, 0s);
    remEqualTestOuter<short, short>(42s, 8s, 2s, -2s, -2s, 2s);
    remEqualTestOuter<short, long>(100s, 26l, 22s, -22s, -22s, 22s);
    // Lhs long
    remEqualTestOuter<long, int>(42l, 7, -0l, -0l, 0l, 0l);
    remEqualTestOuter<long, short>(42l, 10s, 2l, -2l, -2l, 2l);
    remEqualTestOuter<long, long>(10932847123l, 234324l, 226579l, -226579l, -226579l, 226579l);
    // Lhs byte
    remEqualTestInner<byte, byte>(cast<byte>(42), cast<byte>(41), cast<byte>(1));
}

// ------------------------------------------ <<= -----------------------------------------

p shlEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs <<= rhs;
    assert lhs == expectedResult;
}

p shlEqualTest() {
    // Lhs int
    shlEqualTestInner<int, int>(5, 3, 40);
    shlEqualTestInner<int, short>(5, 2s, 20);
    shlEqualTestInner<int, long>(5, 4l, 80);
    // Lhs short
    shlEqualTestInner<short, int>(8s, 2, 32s);
    shlEqualTestInner<short, short>(8s, 1s, 16s);
    shlEqualTestInner<short, long>(8s, 6l, 512s);
    // Lhs long
    shlEqualTestInner<long, int>(7l, 7, 896l);
    shlEqualTestInner<long, short>(7l, 10s, 7168l);
    shlEqualTestInner<long, long>(1234876l, 21l, 2589722673152l);
    // Lhs byte
    shlEqualTestInner<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(84));
}

// ------------------------------------------ >>= -----------------------------------------

p shrEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs >>= rhs;
    assert lhs == expectedResult;
}

p shrEqualTest() {
    // Lhs int
    shrEqualTestInner<int, int>(5, 3, 0);
    shrEqualTestInner<int, short>(5, 2s, 1);
    shrEqualTestInner<int, long>(5, 1l, 2);
    // Lhs short
    shrEqualTestInner<short, int>(8s, 2, 2s);
    shrEqualTestInner<short, short>(8s, 1s, 4s);
    shrEqualTestInner<short, long>(8s, 3l, 1s);
    // Lhs long
    shrEqualTestInner<long, int>(23425l, 7, 183l);
    shrEqualTestInner<long, short>(34587334534l, 10s, 33776693l);
    shrEqualTestInner<long, long>(1234876l, 21l, 0l);
    // Lhs byte
    shrEqualTestInner<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(21));
}

// ------------------------------------------ &= ------------------------------------------

p andEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs &= rhs;
    assert lhs == expectedResult;
}

p andEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    andEqualTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p andEqualTest() {
    // Lhs int
    andEqualTestOuter<int, int>(5, 3, 1);
    andEqualTestOuter<int, short>(5, 2s, 0);
    andEqualTestOuter<int, long>(5, 1l, 1);
    // Lhs short
    andEqualTestOuter<short, int>(8s, 2, 0s);
    andEqualTestOuter<short, short>(8s, 1s, 0s);
    andEqualTestOuter<short, long>(8s, 3l, 0s);
    // Lhs long
    andEqualTestOuter<long, int>(23425l, 7, 1l);
    andEqualTestOuter<long, short>(34587334534l, 10s, 2l);
    andEqualTestOuter<long, long>(1234876l, 21l, 20l);
    // Lhs byte
    andEqualTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(0));
}

// ------------------------------------------ |= ------------------------------------------

p orEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs |= rhs;
    assert lhs == expectedResult;
}

p orEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    orEqualTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p orEqualTest() {
    // Lhs int
    orEqualTestOuter<int, int>(5, 3, 7);
    orEqualTestOuter<int, short>(5, 2s, 7);
    orEqualTestOuter<int, long>(5, 1l, 5);
    // Lhs short
    orEqualTestOuter<short, int>(8s, 2, 10s);
    orEqualTestOuter<short, short>(8s, 1s, 9s);
    orEqualTestOuter<short, long>(8s, 3l, 11s);
    // Lhs long
    orEqualTestOuter<long, int>(23425l, 7, 23431l);
    orEqualTestOuter<long, short>(34587334534l, 10s, 34587334542l);
    orEqualTestOuter<long, long>(1234876l, 21l, 1234877l);
    // Lhs byte
    orEqualTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(43));
}

// ------------------------------------------ ^= ------------------------------------------

p xorEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs ^= rhs;
    assert lhs == expectedResult;
}

p xorEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    xorEqualTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p xorEqualTest() {
    // Lhs int
    xorEqualTestOuter<int, int>(5, 3, 6);
    xorEqualTestOuter<int, short>(5, 2s, 7);
    xorEqualTestOuter<int, long>(5, 1l, 4);
    // Lhs short
    xorEqualTestOuter<short, int>(8s, 2, 10s);
    xorEqualTestOuter<short, short>(8s, 1s, 9s);
    xorEqualTestOuter<short, long>(8s, 3l, 11s);
    // Lhs long
    xorEqualTestOuter<long, int>(23425l, 7, 23430l);
    xorEqualTestOuter<long, short>(34587334534l, 10s, 34587334540l);
    xorEqualTestOuter<long, long>(1234876l, 21l, 1234857l);
    // Lhs byte
    xorEqualTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(43));
}

// ------------------------------------------ ^ ------------------------------------------

p bitwiseXorTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs ^ rhs;
    assert actualResult == expectedResult;
}

p bitwiseXorTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    bitwiseXorTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p bitwiseXorTest() {
    // Lhs int
    bitwiseXorTestOuter<int, int>(5, 3, 6);
    // Lhs short
    bitwiseXorTestOuter<short, short>(8s, 1s, 9s);
    // Lhs long
    bitwiseXorTestOuter<long, long>(1234876l, 21l, 1234857l);
    // Lhs byte
    bitwiseXorTestOuter<byte, byte>(cast<byte>(15), cast<byte>(23), cast<byte>(24));
    // Lhs bool
    bitwiseXorTestOuter<bool, bool>(false, false, false);
    bitwiseXorTestOuter<bool, bool>(false, true, true);
    bitwiseXorTestOuter<bool, bool>(true, false, true);
    bitwiseXorTestOuter<bool, bool>(true, true, false);
}

// ------------------------------------------ | ------------------------------------------

p bitwiseOrTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs | rhs;
    assert actualResult == expectedResult;
}

p bitwiseOrTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    bitwiseOrTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p bitwiseOrTest() {
    // Lhs int
    bitwiseOrTestOuter<int, int>(5, 3, 7);
    // Lhs short
    bitwiseOrTestOuter<short, short>(8s, 1s, 9s);
    // Lhs long
    bitwiseOrTestOuter<long, long>(1234876l, 21l, 1234877l);
    // Lhs byte
    bitwiseOrTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(43));
    // Lhs bool
    bitwiseOrTestOuter<bool, bool>(false, false, false);
    bitwiseOrTestOuter<bool, bool>(false, true, true);
    bitwiseOrTestOuter<bool, bool>(true, false, true);
    bitwiseOrTestOuter<bool, bool>(true, true, true);
}

// ------------------------------------------ & ------------------------------------------

p bitwiseAndTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs & rhs;
    assert actualResult == expectedResult;
}

p bitwiseAndTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    bitwiseAndTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p bitwiseAndTest() {
    // Lhs int
    bitwiseAndTestOuter<int, int>(5, 3, 1);
    // Lhs short
    bitwiseAndTestOuter<short, short>(8s, 1s, 0s);
    // Lhs long
    bitwiseAndTestOuter<long, long>(1234876l, 21l, 20l);
    // Lhs byte
    bitwiseAndTestOuter<byte, byte>(cast<byte>(15), cast<byte>(23), cast<byte>(7));
    // Lhs bool
    bitwiseAndTestOuter<bool, bool>(false, false, false);
    bitwiseAndTestOuter<bool, bool>(false, true, false);
    bitwiseAndTestOuter<bool, bool>(true, false, false);
    bitwiseAndTestOuter<bool, bool>(true, true, true);
}

// ------------------------------------------ == -----------------------------------------

p equalTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs == rhs;
    assert actualResult == expectedResult;
}

p equalTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    equalTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    equalTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    equalTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    equalTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p equalTest() {
    // Lhs is ptr
    int i = 213;
    int* iPtr = &i;
    equalTestInner<int*, int*>(iPtr, iPtr, false);
    equalTestInner<int*, unsigned long>(iPtr, 0ul, false);
    // Lhs double
    equalTestOuter<double, int>(87.0, 87, true, false, false, true);
    equalTestOuter<double, short>(14.0, 14s, true, false, false, true);
    equalTestOuter<double, long>(2349234.0, 2349234l, true, false, false, true);
    // Lhs int
    equalTestOuter<int, double>(12345, 12345.0, true, false, false, true);
    equalTestOuter<int, int>(5, 5, true, false, false, true);
    equalTestOuter<int, short>(-234, -234s, true, false, false, true);
    equalTestOuter<int, long>(-9999999, 9999999l, false, true, true, false);
    equalTestInner<int, char>(67, 'C', true);
    // Lhs short
    equalTestOuter<short, double>(12345s, 12345.0, true, false, false, true);
    equalTestOuter<short, int>(5s, 5, true, false, false, true);
    equalTestOuter<short, short>(-234s, -234s, true, false, false, true);
    equalTestOuter<short, long>(-999s, 999l, false, true, true, false);
    equalTestInner<short, char>(68s, 'D', true);
    // Lhs long
    equalTestOuter<long, double>(12345l, 12345.0, true, false, false, true);
    equalTestOuter<long, int>(5l, 5, true, false, false, true);
    equalTestOuter<long, short>(-234l, -234s, true, false, false, true);
    equalTestOuter<long, long>(-999l, 999l, false, true, true, false);
    equalTestInner<long, char>(68l, 'D', true);
    // Lhs byte
    equalTestInner<byte, byte>(cast<byte>(15), cast<byte>(15), true);
    // Lhs char
    equalTestInner<char, int>('x', -15, false);
    equalTestInner<char, short>('5', 53s, true);
    equalTestInner<char, long>('+', 43l, true);
    equalTestInner<char, char>('#', '#', true);
    // Lhs string
    equalTestInner<string, string>("this is a test", "this is a test", true);
    equalTestInner<string, string>("string", "strong", false);
    String strA = String("this is a test");
    String strB = String("strong");
    equalTestInner<string, string>("this is a test", strA.getRaw(), true);
    equalTestInner<string, string>("string", strB.getRaw(), false);
    // Lhs bool
    equalTestInner<bool, bool>(false, false, false);
    equalTestInner<bool, bool>(false, true, true);
    equalTestInner<bool, bool>(true, false, true);
    equalTestInner<bool, bool>(true, true, false);
    // Lhs function
    const dyn funcA = f<int>(bool _b, double _d) { return 123; };
    const dyn funcB = f<int>(bool _b, double _d) { return 456; };
    equalTestInner<f<int>(bool, double), f<int>(bool, double)>(funcA, funcA, true);
    equalTestInner<f<int>(bool, double), f<int>(bool, double)>(funcA, funcB, false);
    // Lhs procedure
    const dyn procA = p(string _s, char _c) {};
    const dyn procB = p(string _s, char _c) {};
    equalTestInner<p(string, char), p(string, char)>(procA, procA, true);
    equalTestInner<p(string, char), p(string, char)>(procA, procB, false);
}

// ------------------------------------------ != -----------------------------------------

p notEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs != rhs;
    assert actualResult == expectedResult;
}

p notEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    notEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    notEqualTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    notEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    notEqualTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p notEqualTest() {
    // Lhs is ptr
    int i = 213;
    int* iPtr = &i;
    notEqualTestInner<int*, int*>(iPtr, iPtr, true);
    notEqualTestInner<int*, unsigned long>(iPtr, 0ul, false);
    // Lhs double
    notEqualTestOuter<double, int>(87.0, 87, false, true, true, false);
    notEqualTestOuter<double, short>(14.0, 14s, false, true, true, false);
    notEqualTestOuter<double, long>(2349234.0, 2349234l, false, true, true, false);
    // Lhs int
    notEqualTestOuter<int, double>(12345, 12345.0, false, true, true, false);
    notEqualTestOuter<int, int>(5, 5, false, true, true, false);
    notEqualTestOuter<int, short>(-234, -234s, false, true, true, false);
    notEqualTestOuter<int, long>(-9999999, 9999999l, true, false, false, true);
    notEqualTestInner<int, char>(67, 'C', false);
    // Lhs short
    notEqualTestOuter<short, double>(12345s, 12345.0, false, true, true, false);
    notEqualTestOuter<short, int>(5s, 5, false, true, true, false);
    notEqualTestOuter<short, short>(-234s, -234s, false, true, true, false);
    notEqualTestOuter<short, long>(-999s, 999l, true, false, false, true);
    notEqualTestInner<short, char>(68s, 'D', false);
    // Lhs long
    notEqualTestOuter<long, double>(12345l, 12345.0, false, true, true, false);
    notEqualTestOuter<long, int>(5l, 5, false, true, true, false);
    notEqualTestOuter<long, short>(-234l, -234s, false, true, true, false);
    notEqualTestOuter<long, long>(-999l, 999l, true, false, false, true);
    notEqualTestInner<long, char>(68l, 'D', false);
    // Lhs byte
    notEqualTestInner<byte, byte>(cast<byte>(15), cast<byte>(15), false);
    // Lhs char
    notEqualTestInner<char, int>('x', -15, true);
    notEqualTestInner<char, short>('5', 53s, false);
    notEqualTestInner<char, long>('+', 43l, false);
    notEqualTestInner<char, char>('#', '#', false);
    // Lhs string
    notEqualTestInner<string, string>("this is a test", "this is a test", false);
    notEqualTestInner<string, string>("string", "strong", true);
    String strA = String("this is a test");
    String strB = String("strong");
    notEqualTestInner<string, string>("this is a test", strA.getRaw(), false);
    notEqualTestInner<string, string>("string", strB.getRaw(), true);
    // Lhs bool
    notEqualTestInner<bool, bool>(false, false, true);
    notEqualTestInner<bool, bool>(false, true, false);
    notEqualTestInner<bool, bool>(true, false, false);
    notEqualTestInner<bool, bool>(true, true, true);
    // Lhs function
    const dyn funcA = f<int>(bool _b, double _d) { return 123; };
    const dyn funcB = f<int>(bool _b, double _d) { return 456; };
    notEqualTestInner<f<int>(bool, double), f<int>(bool, double)>(funcA, funcA, false);
    notEqualTestInner<f<int>(bool, double), f<int>(bool, double)>(funcA, funcB, true);
    // Lhs procedure
    const dyn procA = p(string _s, char _c) {};
    const dyn procB = p(string _s, char _c) {};
    notEqualTestInner<p(string, char), p(string, char)>(procA, procA, false);
    notEqualTestInner<p(string, char), p(string, char)>(procA, procB, true);
}

// ------------------------------------------ < ------------------------------------------

p lessTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs < rhs;
    assert actualResult == expectedResult;
}

p lessTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    lessTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    lessTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    lessTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    lessTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p lessTest() {
    // Lhs double
    lessTestOuter<double, double>(87.123, 87.124, true, false, false, true);
    lessTestOuter<double, int>(87.0, 88, true, false, false, true);
    lessTestOuter<double, short>(14.0, 15s, true, false, false, true);
    lessTestOuter<double, long>(2349234.0, 2349235l, true, false, false, true);
    // Lhs int
    lessTestOuter<int, double>(12345, 12345.1, true, false, false, true);
    lessTestOuter<int, int>(5, 6, true, false, false, true);
    lessTestOuter<int, short>(-234, -233s, true, false, false, true);
    lessTestOuter<int, long>(9999999, -9999999l, false, true, true, false);
    // Lhs short
    lessTestOuter<short, double>(12345s, 12345.423, true, false, false, true);
    lessTestOuter<short, int>(5s, 6, true, false, false, true);
    lessTestOuter<short, short>(-234s, -233s, true, false, false, true);
    lessTestOuter<short, long>(999s, -999l, false, true, true, false);
    // Lhs long
    lessTestOuter<long, double>(12345l, 12345.1, true, false, false, true);
    lessTestOuter<long, int>(5l, 6, true, false, false, true);
    lessTestOuter<long, short>(-234l, -233s, true, false, false, true);
    lessTestOuter<long, long>(999l, -999l, false, true, true, false);
    // Lhs byte
    lessTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), true);
    // Lhs char
    lessTestInner<char, char>('#', '#', false);
}

// ------------------------------------------ > ------------------------------------------

p greaterTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs > rhs;
    assert actualResult == expectedResult;
}

p greaterTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    greaterTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    greaterTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    greaterTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    greaterTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p greaterTest() {
    // Lhs double
    greaterTestOuter<double, double>(87.123, 87.124, false, true, true, false);
    greaterTestOuter<double, int>(87.0, 88, false, true, true, false);
    greaterTestOuter<double, short>(14.0, 15s, false, true, true, false);
    greaterTestOuter<double, long>(2349234.0, 2349235l, false, true, true, false);
    // Lhs int
    greaterTestOuter<int, double>(12345, 12345.1, false, true, true, false);
    greaterTestOuter<int, int>(5, 6, false, true, true, false);
    greaterTestOuter<int, short>(-234, -233s, false, true, true, false);
    greaterTestOuter<int, long>(9999999, -9999999l, true, false, false, true);
    // Lhs short
    greaterTestOuter<short, double>(12345s, 12345.423, false, true, true, false);
    greaterTestOuter<short, int>(5s, 6, false, true, true, false);
    greaterTestOuter<short, short>(-234s, -233s, false, true, true, false);
    greaterTestOuter<short, long>(999s, -999l, true, false, false, true);
    // Lhs long
    greaterTestOuter<long, double>(12345l, 12345.1, false, true, true, false);
    greaterTestOuter<long, int>(5l, 6, false, true, true, false);
    greaterTestOuter<long, short>(-234l, -233s, false, true, true, false);
    greaterTestOuter<long, long>(999l, -999l, true, false, false, true);
    // Lhs byte
    greaterTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), false);
    // Lhs char
    greaterTestInner<char, char>('#', '#', false);
}

// ------------------------------------------ <= -----------------------------------------

p lessEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs <= rhs;
    assert actualResult == expectedResult;
}

p lessEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    lessEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    lessEqualTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    lessEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    lessEqualTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p lessEqualTest() {
    // Lhs double
    lessEqualTestOuter<double, double>(87.123, 87.124, true, false, false, true);
    lessEqualTestOuter<double, int>(87.0, 88, true, false, false, true);
    lessEqualTestOuter<double, short>(14.0, 15s, true, false, false, true);
    lessEqualTestOuter<double, long>(2349234.0, 2349235l, true, false, false, true);
    // Lhs int
    lessEqualTestOuter<int, double>(12345, 12345.1, true, false, false, true);
    lessEqualTestOuter<int, int>(5, 6, true, false, false, true);
    lessEqualTestOuter<int, short>(-234, -233s, true, false, false, true);
    lessEqualTestOuter<int, long>(9999999, -9999999l, false, true, true, false);
    // Lhs short
    lessEqualTestOuter<short, double>(12345s, 12345.423, true, false, false, true);
    lessEqualTestOuter<short, int>(5s, 6, true, false, false, true);
    lessEqualTestOuter<short, short>(-234s, -233s, true, false, false, true);
    lessEqualTestOuter<short, long>(999s, -999l, false, true, true, false);
    // Lhs long
    lessEqualTestOuter<long, double>(12345l, 12345.1, true, false, false, true);
    lessEqualTestOuter<long, int>(5l, 6, true, false, false, true);
    lessEqualTestOuter<long, short>(-234l, -233s, true, false, false, true);
    lessEqualTestOuter<long, long>(999l, -999l, false, true, true, false);
    // Lhs byte
    lessEqualTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), true);
    // Lhs char
    lessEqualTestInner<char, char>('#', '#', true);
}

// ------------------------------------------ >= -----------------------------------------

p greaterEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs >= rhs;
    assert actualResult == expectedResult;
}

p greaterEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    greaterEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    greaterEqualTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    greaterEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    greaterEqualTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p greaterEqualTest() {
    // Lhs double
    greaterEqualTestOuter<double, double>(87.123, 87.124, false, true, true, false);
    greaterEqualTestOuter<double, int>(87.0, 88, false, true, true, false);
    greaterEqualTestOuter<double, short>(14.0, 15s, false, true, true, false);
    greaterEqualTestOuter<double, long>(2349234.0, 2349235l, false, true, true, false);
    // Lhs int
    greaterEqualTestOuter<int, double>(12345, 12345.1, false, true, true, false);
    greaterEqualTestOuter<int, int>(5, 6, false, true, true, false);
    greaterEqualTestOuter<int, short>(-234, -233s, false, true, true, false);
    greaterEqualTestOuter<int, long>(9999999, -9999999l, true, false, false, true);
    // Lhs short
    greaterEqualTestOuter<short, double>(12345s, 12345.423, false, true, true, false);
    greaterEqualTestOuter<short, int>(5s, 6, false, true, true, false);
    greaterEqualTestOuter<short, short>(-234s, -233s, false, true, true, false);
    greaterEqualTestOuter<short, long>(999s, -999l, true, false, false, true);
    // Lhs long
    greaterEqualTestOuter<long, double>(12345l, 12345.1, false, true, true, false);
    greaterEqualTestOuter<long, int>(5l, 6, false, true, true, false);
    greaterEqualTestOuter<long, short>(-234l, -233s, false, true, true, false);
    greaterEqualTestOuter<long, long>(999l, -999l, true, false, false, true);
    // Lhs byte
    greaterEqualTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), false);
    // Lhs char
    greaterEqualTestInner<char, char>('#', '#', true);
}

// ------------------------------------------ << -----------------------------------------

p shlTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs << rhs;
    assert actualResult == expectedResult;
}

p shlTest() {
    // Lhs int
    shlTestInner<int, int>(5, 3, 40);
    shlTestInner<int, short>(5, 2s, 20);
    shlTestInner<int, long>(5, 4l, 80);
    // Lhs short
    shlTestInner<short, int>(8s, 2, 32s);
    shlTestInner<short, short>(8s, 1s, 16s);
    shlTestInner<short, long>(8s, 6l, 512s);
    // Lhs long
    shlTestInner<long, int>(7l, 7, 896l);
    shlTestInner<long, short>(7l, 10s, 7168l);
    shlTestInner<long, long>(1234876l, 21l, 2589722673152l);
    // Lhs byte
    shlTestInner<byte, int>(cast<byte>(3), 2, cast<byte>(12));
    shlTestInner<byte, short>(cast<byte>(3), 2s, cast<byte>(12));
    shlTestInner<byte, long>(cast<byte>(3), 2l, cast<byte>(12));
    shlTestInner<byte, byte>(cast<byte>(3), cast<byte>(2), cast<byte>(12));
}

// ------------------------------------------ >> -----------------------------------------

p shrTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs >> rhs;
    assert actualResult == expectedResult;
}

p shrTest() {
    // Lhs int
    shrTestInner<int, int>(5, 3, 0);
    shrTestInner<int, short>(5, 2s, 1);
    shrTestInner<int, long>(5, 1l, 2);
    // Lhs short
    shrTestInner<short, int>(8s, 2, 2s);
    shrTestInner<short, short>(8s, 1s, 4s);
    shrTestInner<short, long>(8s, 3l, 1s);
    // Lhs long
    shrTestInner<long, int>(23425l, 7, 183l);
    shrTestInner<long, short>(34587334534l, 10s, 33776693l);
    shrTestInner<long, long>(1234876l, 21l, 0l);
    // Lhs byte
    shrTestInner<byte, int>(cast<byte>(12), 2, cast<byte>(3));
    shrTestInner<byte, short>(cast<byte>(12), 2s, cast<byte>(3));
    shrTestInner<byte, long>(cast<byte>(12), 2l, cast<byte>(3));
    shrTestInner<byte, byte>(cast<byte>(12), cast<byte>(2), cast<byte>(3));
}

// ------------------------------------------ + -------------------------------------------

p plusTestInner<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult) {
    const TRes actualResult = lhs + rhs;
    assert actualResult == expectedResult;
}

p plusTestInnerUnsafe<TRhs>(int* lhs, const TRhs rhs, const int* expectedResult) {
    unsafe {
        const int* actualResult = lhs + rhs;
        assert actualResult == expectedResult;
    }
}

p plusTestOuter<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult1, const TRes expectedResult2, const TRes expectedResult3, const TRes expectedResult4) {
    plusTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    plusTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    plusTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    plusTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p plusTest() {
    // Lhs is double
    plusTestOuter<double, double, double>(1.234, 98.7654, 99.9994, -99.9994, 97.5314, -97.5314);
    plusTestOuter<double, int, double>(1.234, 98, 99.234, -99.234, 96.766, -96.766);
    plusTestOuter<double, short, double>(1.234, 98s, 99.234, -99.234, 96.766, -96.766);
    plusTestOuter<double, long, double>(1.234, 98l, 99.234, -99.234, 96.766, -96.766);
    // Lhs is int
    plusTestOuter<int, double, double>(78, 674.45, 752.45, -752.45, 596.45, -596.45);
    plusTestOuter<int, int, int>(78, 674, 752, -752, 596, -596);
    plusTestOuter<int, short, int>(78, 7s, 85, -85, -71, 71);
    plusTestOuter<int, long, long>(78, 2384723l, 2384801l, -2384801l, 2384645l, -2384645l);
    // Lhs is short
    plusTestOuter<short, double, double>(78s, 674.76, 752.76, -752.76, 596.76, -596.76);
    plusTestOuter<short, int, int>(78s, 674, 752, -752, 596, -596);
    plusTestOuter<short, short, short>(78s, 7s, 85s, -85s, -71s, 71s);
    plusTestOuter<short, long, long>(78s, 2384723l, 2384801l, -2384801l, 2384645l, -2384645l);
    // Lhs is long
    plusTestOuter<long, double, double>(78l, 674.91, 752.91, -752.91, 596.91, -596.91);
    plusTestOuter<long, int, long>(78l, 674, 752l, -752l, 596l, -596l);
    plusTestOuter<long, short, long>(78l, 7s, 85l, -85l, -71l, 71l);
    plusTestOuter<long, long, long>(78l, 2384723l, 2384801l, -2384801l, 2384645l, -2384645l);
    // Lhs is byte
    plusTestInner<byte, byte, byte>(cast<byte>(5), cast<byte>(6), cast<byte>(11));
    // Lhs is ptr
    int[5] input = [0, 0, 0, 0, 0];
    plusTestInnerUnsafe(&input[2], 2, &input[4]);
    plusTestInnerUnsafe(&input[2], -2, &input[0]);
    plusTestInnerUnsafe(&input[2], 2s, &input[4]);
    plusTestInnerUnsafe(&input[2], -2s, &input[0]);
    plusTestInnerUnsafe(&input[2], 2l, &input[4]);
    plusTestInnerUnsafe(&input[2], -2l, &input[0]);
}

// ------------------------------------------ - -------------------------------------------

p minusTestInner<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult) {
    const TRes actualResult = lhs - rhs;
    assert actualResult == expectedResult;
}

p minusTestInnerUnsafe<TRhs>(int* lhs, const TRhs rhs, const int* expectedResult) {
    unsafe {
        const int* actualResult = lhs - rhs;
        assert actualResult == expectedResult;
    }
}

p minusTestOuter<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult1, const TRes expectedResult2, const TRes expectedResult3, const TRes expectedResult4) {
    minusTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    minusTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    minusTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    minusTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p minusTest() {
    // Lhs is double
    minusTestOuter<double, double, double>(1.234, 98.7654, -97.5314, 97.5314, -99.9994, 99.9994);
    minusTestOuter<double, int, double>(1.234, 98, -96.766, 96.766, -99.234, 99.234);
    minusTestOuter<double, short, double>(1.234, 98s, -96.766, 96.766, -99.234, 99.234);
    minusTestOuter<double, long, double>(1.234, 98l, -96.766, 96.766, -99.234, 99.234);
    // Lhs is int
    minusTestOuter<int, double, double>(78, 674.45, -596.45, 596.45, -752.45, 752.45);
    minusTestOuter<int, int, int>(78, 674, -596, 596, -752, 752);
    minusTestOuter<int, short, int>(78, 7s, 71, -71, -85, 85);
    minusTestOuter<int, long, long>(78, 2384723l, -2384645l, 2384645l, -2384801l, 2384801l);
    // Lhs is short
    minusTestOuter<short, double, double>(78s, 674.76, -596.76, 596.76, -752.76, 752.76);
    minusTestOuter<short, int, int>(78s, 674, -596, 596, -752, 752);
    minusTestOuter<short, short, short>(78s, 7s, 71s, -71s, -85s, 85s);
    minusTestOuter<short, long, long>(78s, 2384723l, -2384645l, 2384645l, -2384801l, 2384801l);
    // Lhs is long
    minusTestOuter<long, double, double>(78l, 674.91, -596.91, 596.91, -752.91, 752.91);
    minusTestOuter<long, int, long>(78l, 674, -596l, 596l, -752l, 752l);
    minusTestOuter<long, short, long>(78l, 7s, 71l, -71l, -85l, 85l);
    minusTestOuter<long, long, long>(78l, 2384723l, -2384645l, 2384645l, -2384801l, 2384801l);
    // Lhs is byte
    minusTestInner<byte, byte, byte>(cast<byte>(6), cast<byte>(5), cast<byte>(1));
    // Lhs is ptr
    int[5] input = [0, 0, 0, 0, 0];
    minusTestInnerUnsafe(&input[2], 2, &input[0]);
    minusTestInnerUnsafe(&input[2], -2, &input[4]);
    minusTestInnerUnsafe(&input[2], 2s, &input[0]);
    minusTestInnerUnsafe(&input[2], -2s, &input[4]);
    minusTestInnerUnsafe(&input[2], 2l, &input[0]);
    minusTestInnerUnsafe(&input[2], -2l, &input[4]);
}

// ------------------------------------------ * -------------------------------------------

p mulTestInner<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult) {
    const TRes actualResult = lhs * rhs;
    assert actualResult == expectedResult;
}

p mulTestOuter<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult1, const TRes expectedResult2, const TRes expectedResult3, const TRes expectedResult4) {
    mulTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    mulTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    mulTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    mulTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p mulTest() {
    // Lhs is double
    mulTestOuter<double, double, double>(1.23, 98.76, 121.4748, 121.4748, -121.4748, -121.4748);
    mulTestOuter<double, int, double>(1.234, 98, 120.932, 120.932, -120.932, -120.932);
    mulTestOuter<double, short, double>(1.234, 98s, 120.932, 120.932, -120.932, -120.932);
    mulTestOuter<double, long, double>(1.234, 98l, 120.932, 120.932, -120.932, -120.932);
    // Lhs is int
    mulTestOuter<int, double, double>(78, 674.4, 52603.2, 52603.2, -52603.2, -52603.2);
    mulTestOuter<int, int, int>(78, 674, 52572, 52572, -52572, -52572);
    mulTestOuter<int, short, int>(78, 7s, 546, 546, -546, -546);
    mulTestOuter<int, long, long>(78, 2384723l, 186008394l, 186008394l, -186008394l, -186008394l);
    // Lhs is short
    mulTestOuter<short, double, double>(78s, 674.76, 52631.28, 52631.28, -52631.28, -52631.28);
    mulTestOuter<short, int, int>(78s, 674, 52572, 52572, -52572, -52572);
    mulTestOuter<short, short, short>(78s, 7s, 546s, 546s, -546s, -546s);
    mulTestOuter<short, long, long>(78s, 2384723l, 186008394l, 186008394l, -186008394l, -186008394l);
    // Lhs is long
    mulTestOuter<long, double, double>(78l, 674.9, 52642.2, 52642.2, -52642.2, -52642.2);
    mulTestOuter<long, int, long>(78l, 674, 52572l, 52572l, -52572l, -52572l);
    mulTestOuter<long, short, long>(78l, 7s, 546l, 546l, -546l, -546l);
    mulTestOuter<long, long, long>(78l, 2384723l, 186008394l, 186008394l, -186008394l, -186008394l);
    // Lhs is byte
    mulTestInner<byte, byte, byte>(cast<byte>(6), cast<byte>(5), cast<byte>(30));
}

// ------------------------------------------ / -------------------------------------------

p divTestInner<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult) {
    const TRes actualResult = lhs / rhs;
    assert actualResult == expectedResult;
}

p divTestOuter<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult1, const TRes expectedResult2, const TRes expectedResult3, const TRes expectedResult4) {
    divTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    divTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    divTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    divTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p divTest() {
    // Lhs is double
    divTestOuter<double, double, double>(121.4748, 98.76, 1.23, 1.23, -1.23, -1.23);
    divTestOuter<double, int, double>(120.932, 98, 1.234, 1.234, -1.234, -1.234);
    divTestOuter<double, short, double>(120.932, 98s, 1.234, 1.234, -1.234, -1.234);
    divTestOuter<double, long, double>(120.932, 98l, 1.234, 1.234, -1.234, -1.234);
    // Lhs is int
    divTestOuter<int, double, double>(500, 50.0, 10.0, 10.0, -10.0, -10.0);
    divTestOuter<int, int, int>(52572, 674, 78, 78, -78, -78);
    divTestOuter<int, short, int>(546, 7s, 78, 78, -78, -78);
    divTestOuter<int, long, long>(186008394, 2384723l, 78l, 78l, -78l, -78l);
    // Lhs is short
    divTestOuter<short, double, double>(6s, 1.5, 4.0, 4.0, -4.0, -4.0);
    divTestOuter<short, int, int>(10s, 5, 2, 2, -2, -2);
    divTestOuter<short, short, short>(546s, 7s, 78s, 78s, -78s, -78s);
    divTestOuter<short, long, long>(78s, 2384723l, 0l, 0l, -0l, -0l);
    // Lhs is long
    divTestOuter<long, double, double>(52642l, 2.5, 21056.8, 21056.8, -21056.8, -21056.8);
    divTestOuter<long, int, long>(52572l, 674, 78l, 78l, -78l, -78l);
    divTestOuter<long, short, long>(546l, 7s, 78l, 78l, -78l, -78l);
    divTestOuter<long, long, long>(186008394l, 2384723l, 78l, 78l, -78l, -78l);
    // Lhs is byte
    divTestInner<byte, byte, byte>(cast<byte>(30), cast<byte>(5), cast<byte>(6));
}

// ------------------------------------------ % -------------------------------------------

p remTestInner<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult) {
    const TRes actualResult = lhs % rhs;
    //printf("actualResult: %d, expectedResult: %d\n", actualResult, expectedResult);
    //printf("actualResult: %f, expectedResult: %f\n", actualResult, expectedResult);
    assert actualResult == expectedResult;
}

p remTestOuter<TLhs, TRhs, TRes>(TLhs lhs, const TRhs rhs, const TRes expectedResult1, const TRes expectedResult2, const TRes expectedResult3, const TRes expectedResult4) {
    remTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    remTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    remTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    remTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p remTest() {
    // Lhs is double
    remTestOuter<double, double, double>(121.0, 5.5, 0.0, -0.0, -0.0, 0.0);
    // Lhs is int
    remTestOuter<int, int, int>(52572, 674, 0, 0, -0, -0);
    remTestOuter<int, short, int>(546, 8s, 2, -2, -2, 2);
    remTestOuter<int, long, long>(186008394, 238l, 208l, -208l, -208l, 208l);
    // Lhs is short
    remTestOuter<short, int, int>(10s, 5, 0, -0, -0, 0);
    remTestOuter<short, short, short>(546s, 9s, 6s, -6s, -6s, 6s);
    remTestOuter<short, long, long>(78s, 78l, 0l, -0l, -0l, 0l);
    // Lhs is long
    remTestOuter<long, int, long>(52572l, 1, 0l, -0l, -0l, 0l);
    remTestOuter<long, short, long>(546l, 11s, 7l, -7l, -7l, 7l);
    remTestOuter<long, long, long>(186008394l, 186008393l, 1l, -1l, -1l, 1l);
}

f<int> main() {
    plusEqualTest();    // x += y
    minusEqualTest();   // x -= y
    mulEqualTest();     // x *= y
    divEqualTest();     // x /= y
    remEqualTest();     // x %= y
    shlEqualTest();     // x <<= y
    shrEqualTest();     // x >>= y
    andEqualTest();     // x &= y
    orEqualTest();      // x |= y
    xorEqualTest();     // x ^= y
    bitwiseOrTest();    // x | y
    bitwiseXorTest();   // x ^ y
    bitwiseAndTest();   // x & y
    equalTest();        // x == y
    notEqualTest();     // x != y
    lessTest();         // x < y
    greaterTest();      // x > y
    lessEqualTest();    // x <= y
    greaterEqualTest(); // x >= y
    shlTest();          // x << y
    shrTest();          // x >> y
    plusTest();         // x + y
    minusTest();        // x - y
    mulTest();          // x * y
    divTest();          // x / y
    remTest();          // x % y
    printf("All assertions passed!");
}