// Imports
import "std/io/file" as file;

public type Reader struct {
    File inputFile
    char curChar
    char nextChar
    bool metEof
    unsigned long line
    unsigned long col
}

public p Reader.ctor(const string inputFileName) {
    this.inputFile = file.openFile(inputFileName, file::MODE_READ);
    this.cursorPos = 0;
    this.metEof = false;
    this.line = 1;
    this.col = 0;
    // Fill
}

public f<char> Reader.getCurChar() {
    return this.curChar;
}

public f<bool> Reader.expectChar(char expected) {
    bool gotExpected = expected == this.nextChar;
    this.advance();
    return gotExpected;
}

public p Reader.advance() {
    int readChar = this.inputFile.readChar();
    if readChar == -1 {
        metEof = true;
        return;
    }
    this.curChar = this.nextChar;
    this.nextChar = (char) readChar;
}