f<int> main() {
    printf("Output: %s", test);
}