f<int> main() {
    int[7] intArray = { 1, 5, 4, 0, 12, 12345, 9 };
    /*foreach (int index = 2, int item : intArray) {
        printf("Item for index %d, %d\n", index, item);
    }*/
    foreach const int item : intArray {
        printf("Index: %d", idx);
        printf("Item: %d", item);
    }
    /*for dyn i = 1; i < 5; i += 2 {
        printf("Item for index %d, %d", i, intArray[i]);
    }*/
}