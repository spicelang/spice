f<int> main() {
    const unsigned signed int test = 1;
}