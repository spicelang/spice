//import "std/os/os" as os;

// File permission modes
public const int MODE_ALL_RWX   = 0o0000777;
public const int MODE_ALL_RW    = 0o0000666;
public const int MODE_ALL_R     = 0o0000444;

public const int MODE_OWNER_RWX = 0o0000700;
public const int MODE_OWNER_R   = 0o0000400;
public const int MODE_OWNER_W   = 0o0000200;
public const int MODE_OWNER_X   = 0o0000100;

public const int MODE_GROUP_RWX = 0o0000070;
public const int MODE_GROUP_R   = 0o0000040;
public const int MODE_GROUP_W   = 0o0000020;
public const int MODE_GROUP_X   = 0o0000010;

public const int MODE_OTHER_RWX = 0o0000007;
public const int MODE_OTHER_R   = 0o0000004;
public const int MODE_OTHER_W   = 0o0000002;
public const int MODE_OTHER_X   = 0o0000001;

const int F_OK = 0; // File existence
const int X_OK = 1; // Can execute
const int W_OK = 2; // Can write
const int R_OK = 4; // Can read

const int IF_MT  = 0o0170000;
const int IF_DIR = 0o0040000;

type FileStat struct {         // Total size: 46 bytes
    unsigned long st_dev       // ID of the device containing file
    unsigned long st_ino       // Inode number
    long st_nlink              // Number of hard links
    unsigned int st_mode       // File type and mode
    int st_uid                 // User ID of owner
    int st_gid                 // Group ID of owner
    unsigned long st_rdev      // Device ID (if special file)
    long st_size               // Total size in bytes
    long st_blksize            // Block size for filesystem I/O
    long st_blocks             // Number of 512B blocks allocated
    long st_atime              // Time of last access
    unsigned long st_atimensec // Nsecs of last access
    long st_mtime              // Time of last modification
    unsigned long st_mtimensec // Nsecs of last modification
    long st_ctime              // Time of last status change
    unsigned long st_ctimensec // Nsecs of last status change
    long[3] __glibc_reserved0
    int __glibc_reserved1
}

type DirEntry struct {
    unsigned long dInodeNo
    long dOffset
    unsigned short dRecordLen
    char dType
    char* dName
}

type DirStream struct {
    int fileDescriptor

}

// Link external functions
ext<int> mkdir(string, int);
ext<int> rmdir(string);
ext<int> rename(string, string);
ext<int> access(string, int);
ext<int> stat(string, FileStat*);
ext<DirStream*> opendir(string);
ext<int> closedir(DirStream*);
ext<DirEntry*> readdir(DirStream*);

/**
 * Creates an empty directory at the specified path, with the specified mode.
 * Creates at max one directory. If the second last path element does not exist, the operation fails
 *
 * There are predefined constants for the mode available:
 * MODE_ALL_RWX, MODE_ALL_RW, MODE_ALL_R,
 * MODE_OWNER_RWX, MODE_OWNER_R, MODE_OWNER_W, MODE_OWNER_X,
 * MODE_GROUP_RWX, MODE_GROUP_R, MODE_GROUP_W, MODE_GROUP_X,
 * MODE_OTHER_RWX, MODE_OTHER_R, MODE_OTHER_W, MODE_OTHER_X
 *
 * @return Result code of the create operation: 0 = successful, -1 = failed
 */
public f<int> mkDir(string path, int mode) {
    return mkdir(path, mode);
}

/**
 * Creates an empty directory at the specified path, with the specified mode.
 * Unlike mkDir, mkDirs can also create nested path structures.
 *
 * There are predefined constants for the mode available:
 * MODE_ALL_RWX, MODE_ALL_RW, MODE_ALL_R,
 * MODE_OWNER_RWX, MODE_OWNER_R, MODE_OWNER_W, MODE_OWNER_X,
 * MODE_GROUP_RWX, MODE_GROUP_R, MODE_GROUP_W, MODE_GROUP_X,
 * MODE_OTHER_RWX, MODE_OTHER_R, MODE_OTHER_W, MODE_OTHER_X
 *
 * @return Result code of the create operation: 0 = successful, -1 = failed
 */
public f<int> mkDirs(string path, int mode) {
    // ToDo: Implement

    /*char[] pathChars = (char[]) path;
    for int i = 0; i < path.length(); i++ {

    }*/
    return -1;
}

/**
 * Deletes an empty directory at the specified path.
 *
 * @return Result code of the delete operation: 0 = successful, -1 = failed
 */
public f<int> rmDir(string path) {
    return rmdir(path);
}

/**
 * Renames a directory.
 *
 * @return Result code of the rename operation: 0 = successful, -1 = failed
 */
public f<int> renameDir(string oldPath, string newPath) {
    return rename(oldPath, newPath);
}

/**
 * Checks if a directory is existing.
 *
 * @return Existing or not
 */
public f<bool> dirExists(string path) {
    // Check if there exists something, a file or a dir
    if access(path, F_OK) == 0 {
        // Check if it is a dir
        dyn fs = FileStat{};
        if stat(path, &fs) != 0 {
            return false;
        }
        return ((int) fs.st_mode & IF_MT) == IF_DIR;
    }
    return false;
}

/**
 * Lists all files/subdirectories at a given path.
 */
/*public p listDir(string path) {
    // Open the directory stream
    DirStream* dirStream = opendir(path);

    // Return empty array if stream result is nil
    if (dirStream == nil<DirStream*>) { return; }

    dyn dirEntry = &DirEntry{};
    while (dirEntry = readdir(dirStream)) != nil<DirEntry*> {
        printf("Filename: %s\n", dirEntry.dName);
    }
    closedir(dirStream);
}*/