f<int> test(string input) {
    return 12;
}

f<int> main() {
    const f<int>(string) testFct = test;
    int i = testFct();
    printf("Result: %d", i);
}