f<int> main() {
    string test;
    bool b = false;
    if (b) {
        int test = 12;
        printf("%d", test);
    }
    printf("%s", test);
}