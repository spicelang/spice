import "bootstrap/symboltablebuilder/type-chain";

f<int> main() {

}