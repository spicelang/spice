import "std/io/logging";
import "std/io/file";
import "std/io/filepath";

f<int> main() {
     {
        LogFile logFile = LogFile(FilePath("log.txt"), false);
        logFile.logDebug("This is a debug message");
        logFile.logInfo("This is a info message");
        logFile.logWarning("This is a warning message");
        logFile.logError("This is a error message");
    }

    assert fileExists("log.txt");
    Result<String> fileContent = readFile("log.txt");
    String fileText = fileContent.unwrap();
    assert fileText.contains("[debug] This is a debug message");
    assert fileText.contains("[info] This is a info message");
    assert fileText.contains("[warning] This is a warning message");
    assert fileText.contains("[error] This is a error message");
    bool _ = deleteFile("log.txt");
}