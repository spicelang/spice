const int MAX_PATH = 260; // Maximum path length on Windows

ext f<string> GetTempPathA(int, char[]);

public f<string> getTempDir() {
    char[MAX_PATH] path;
    return GetTempPathA(MAX_PATH, path);
}
