const int count;

f<int> main() {
    printf("Test");
}