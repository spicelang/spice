import "std/data/vector";

f<int> main() {

}