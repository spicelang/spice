import "source3" as s3;

public f<int> dummy() {
    return 2 + s3::dummy() + dummy();
}