f<int> main() {
    assert "Test";
    printf("Unreachable");
}