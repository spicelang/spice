type T dyn;
type U dyn;

p printDyn<T>(T a1, U a2) {
    printf("%d", a1 + a2);
}

f<int> main() {
    printDyn<double, int>(1.3, 4);
}