f<int> main() {
    String str = String();
    unsigned long i = 123l;
    str.reserve(i);
}