import "std/data/queue";

f<Queue<String>> getStringQueue() {
    Queue<String> queue;
    queue.push(String("Hello"));
    queue.push(String("World"));
    return queue;
}

f<int> main() {
    const Queue<String> args = getStringQueue();
    foreach unsigned long i, const String& arg : args {
        printf("Arg %d: %s\n", i, arg);
    }
}