type T int|dyn|double;

p foo<T>(T _t) {}

f<int> main() {
    foo(1);
    foo(1.0);
    foo("test");
}