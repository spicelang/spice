type T dyn;

type Optional<T> struct {
    T value
}

p Optional.ctor() {}

f<int> main() {
     dyn oi = Optional();
}