f<int> main1() {
    int i = 0;
    while i < 10 {
        i += 1;
        printf("i is now at: %d\n", i);
    }
}