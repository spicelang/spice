// Std imports

// Own imports

public type Generator struct {

}