// Std imports
import "std/data/vector";
import "std/text/stringstream";

// Own imports
import "bootstrap/source-file-intf";
import "bootstrap/bindings/llvm/llvm" as llvm;

const string SPICE_VERSION = "0.22.5";
const string SPICE_TARGET_OS = "linux";
const string SPICE_TARGET_ARCH = "amd64";
const string SPICE_GIT_HASH = "45fa32083223a49e07259661d3a7130326bb0bfe";
const string SPICE_BUILT_BY = "GitHub Actions";

/**
 * Split the given haystack by the needle and return the last fragment
 *
 * @param haystack Input string
 * @param needle String to search
 * @return Last fragment
 */
public f<String> getLastFragment(const String &haystack, const string needle) {
    const unsigned long index = haystack.rfind(needle);
    return index != -1l ? haystack.getSubstring(index + getRawLength(needle)) : haystack;
}

/**
 * Generate a circular import message from the given source files
 *
 * @param sourceFiles Source files building the circular dependency chain
 * @return Error message
 */
public f<String> getCircularImportMessage(const Vector<const ISourceFile*>& sourceFiles) {
    StringStream message;
    message << "*-----*" << endl();
    message << "|     |" << endl();
    for unsigned long i = 0l; i < sourceFiles.getSize(); i++ {
        const ISourceFile* sourceFile = sourceFiles.get(i);
        if i != 0 { message << "|     |" << endl(); }
        message << "|  ";
        message << sourceFile.getFileName();
        message << endl();
    }
    message << "|     |" << endl();
    message << "*-----*" << endl();
    return message.str();
}

/**
 * Generate the version info string for the Spice driver
 *
 * @return Version info string
 */
public f<String> buildVersionInfo() {
    StringStream versionString;
    versionString << "Spice version: " << SPICE_VERSION << " " << SPICE_TARGET_OS << "/" << SPICE_TARGET_ARCH << endl();
    versionString << "Git hash:      " << SPICE_GIT_HASH << endl();
    versionString << "LLVM version:  " << llvm::getVersionString() << endl();
    versionString << "built by:      " << SPICE_BUILT_BY << endl() << endl();
    versionString << "(c) Marc Auberer 2021-2026";
    String str = versionString.str();
    return str;
}