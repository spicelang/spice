public const int SIZE = 32;
public const int MIN_VALUE = -2147483648;
public const int MAX_VALUE = 2147483647;

const int nSmall = 100;
const string smallsString10 = "0123456789";
const string smallsString100 = "00010203040506070809101112131415161718192021222324252627282930313233343536373839404142434445464748495051525354555657585960616263646566676869707172737475767778798081828384858687888990919293949596979899";

// Converts an int to a double
public f<double> toDouble(int input) {
    // ToDo: Implement
    return 0.0;
}

// Converts an int to a short
public f<short> toShort(int input) {
    return (short) input;
}

// Converts an int to a long
public f<long> toLong(int input) {
    return (long) input;
}

// Converts an int to a byte
public f<byte> toByte(int input) {
    return (byte) input;
}

// Converts an int to a char
public f<char> toChar(int input) {
    return (char) input;
}

// Converts an int to a string
public f<string> toString(int input) {
    // ToDo: Implement (See https://github.com/golang/go/blob/master/src/strconv/itoa.go)
    return "";
}

// Converts an int to a boolean
public f<bool> toBool(int input) {
    return input >= 1;
}

// Helper function: returns the string of a small number
f<string> small(int i) {
    if i < 10 {
        return smallsString10.substring(i, i+1);
    }
    return smallsString100.substring(i*2, i*2+2);
}