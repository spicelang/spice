// TEST: --disable-verifier

f<int> main() {
    printf("Hello World!");
}