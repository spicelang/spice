f<int> main() {
    short arraySize = 6s;
    int[arraySize] array;
    array[2] = 11;
    printf("Item: %d\n", array[0]);
    printf("Item: %d\n", array[1]);
    printf("Item: %d\n", array[2]);
    printf("Item: %d\n", array[3]);
    printf("Item: %d\n", array[4]);
    printf("Item: %d\n", array[5]);
}