const f<int> test(const int& i) {
    printf("%d", i);
}

f<int> main() {
    test(3);
}