import "std/os/dir" as dir;

f<int> main() {
    string path = "./test";
    int r1 = dir.mkDir(path, dir.MODE_ALL_RWX);
    printf("R1: %d\n", r1);
    int r2 = dir.rmDir(path);
    printf("R2: %d\n", r2);
}