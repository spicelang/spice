// Imports
import "../reader/code-loc";

// Enums
public type TokenType enum {
    INVALID = 0,
    // Keyword tokens
    TYPE_DOUBLE = 1,
    TYPE_INT = 2,
    TYPE_SHORT = 3,
    TYPE_LONG = 4,
    TYPE_BYTE = 5,
    TYPE_CHAR = 6,
    TYPE_STRING = 7,
    TYPE_BOOL = 8,
    TYPE_DYN = 9,
    CONST = 10,
    SIGNED = 11,
    UNSIGNED = 12,
    INLINE = 13,
    PUBLIC = 14,
    HEAP = 15,
    COMPOSE = 16,
    F = 17,
    P = 18,
    IF = 19,
    ELSE = 20,
    ASSERT = 21,
    FOR = 22,
    FOREACH = 23,
    DO = 24,
    WHILE = 25,
    IMPORT = 26,
    BREAK = 27,
    CONTINUE = 28,
    RETURN = 29,
    AS = 30,
    STRUCT = 31,
    INTERFACE = 32,
    TYPE = 33,
    ENUM = 34,
    OPERATOR = 35,
    ALIAS = 36,
    UNSAFE = 37,
    NIL = 38,
    MAIN = 39,
    PRINTF = 40,
    SIZEOF = 41,
    ALIGNOF = 42,
    LEN = 43,
    PANIC = 44,
    EXT = 45,
    TRUE = 46,
    FALSE = 47,
    // Operator tokens
    LBRACE = 48,
    RBRACE = 49,
    LPAREN = 50,
    RPAREN = 51,
    LBRACKET = 52,
    RBRACKET = 53,
    LOGICAL_OR = 54,
    LOGICAL_AND = 55,
    BITWISE_OR = 56,
    BITWISE_XOR = 57,
    BITWISE_AND = 58,
    PLUS_PLUS = 59,
    MINUS_MINUS = 60,
    PLUS_EQUAL = 61,
    MINUS_EQUAL = 62,
    MUL_EQUAL = 63,
    DIV_EQUAL = 64,
    REM_EQUAL = 65,
    SHL_EQUAL = 66,
    SHR_EQUAL = 67,
    AND_EQUAL = 68,
    OR_EQUAL = 69,
    XOR_EQUAL = 70,
    PLUS = 71,
    MINUS = 72,
    MUL = 73,
    DIV = 74,
    REM = 75,
    NOT = 76,
    BITWISE_NOT = 77,
    GREATER = 78,
    LESS = 79,
    GREATER_EQUAL = 80,
    LESS_EQUAL = 81,
    SHL = 82,
    SHR = 83,
    EQUAL = 84,
    NOT_EQUAL = 85,
    ASSIGN = 86,
    QUESTION_MARK = 87,
    SEMICOLON = 88,
    COLON = 89,
    COMMA = 90,
    DOT = 91,
    ARROW = 92,
    SCOPE_ACCESS = 93,
    ELLIPSIS = 94,
    FCT_ATTR_PREAMBLE = 95,
    MOD_ATTR_PREAMBLE = 96,
    // Regex tokens
    DOUBLE_LIT = 97,
    INT_LIT = 98,
    SHORT_LIT = 99,
    LONG_LIT = 100,
    CHAR_LIT = 101,
    STRING_LIT = 102,
    IDENTIFIER = 103,
    TYPE_IDENTIFIER = 104,
    // Skipped tokens
    DOC_COMMENT = 105,
    BLOCK_COMMENT = 106,
    LINE_COMMENT = 107,
    EOF = 108
}

public type Token struct {
    public TokenType tokenType
    public String text
    public CodeLoc codeLoc
}

public p Token.ctor(TokenType tokenType) {
    this.tokenType = tokenType;
}

public p Token.ctor(TokenType tokenType, String text, const CodeLoc& codeLoc) {
    this.tokenType = tokenType;
    this.text = text;
    this.codeLoc = codeLoc;
}

public p Token.ctor(TokenType tokenType, string text, const CodeLoc& codeLoc) {
    this.ctor(tokenType, String(text), codeLoc);
}

public p Token.print() {
    printf("Token(type=%d, text=%s, codeLoc=%s)", this.tokenType, this.text, this.codeLoc);
}