public f<bool> isTrue() {
    return true;
}