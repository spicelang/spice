// Link external functions
ext f<heap byte*> malloc(long);
ext p free(heap byte*);

// Add generic type definitions
type T dyn;

/**
 * Node of a DoublyLinkedList
 */
public type Node<T> struct {
    heap Node<T>* prev
    T value
    heap Node<T>* next
}

/**
 * A doubly linked list is a common, dynamically resizable data structure to store uniform data in order.
 * It is characterized by the pointer for every item, pointing to the next one and the pointer, pointing
 * to the previous one.
 */
public type DoublyLinkedList<T> struct {
    heap Node<T>* head
    heap Node<T>* tail
}

public p Node.dtor() {
    if this.next != nil<heap Node<T>*> {
        this.next.dtor();
        free((heap byte*) this.next);
    }
}

public p DoublyLinkedList.insert<T>(T newValue, Node<T>* prevNode = nil<Node<T>*>) {
    // Create new node
    heap Node<T>* newNode;
    unsafe {
        newNode = (heap Node<T>*) malloc(sizeof(type Node<T>) / 8);
    }
    newNode.value = newValue;

    if prevNode != nil<heap Node<T>*> { // Previous node was passed -> insert after this node
        // Link the previous to this one
        newNode.prev = prevNode;
        // Link the next node to this one
        newNode.next = prevNode.next;
        // Link this node to the next node
        prevNode.next.prev = newNode;
        // Link this node to the previous node
        prevNode.next = newNode;

        // Check if the previous node was the last node
        if prevNode == tail {
            this.tail = newNode;
        }
    } else { // No previous node was passed -> insert at head
        newNode.next = this.head;
        this.head = newNode;
    }
}

public p DoublyLinkedList.insertHead<T>(T newValue) {
    this.insert(newValue);
}

public inline p DoublyLinkedList.insertTail<T>(T newValue) {
    this.insert(newValue, this.tail);
}

/*public f<heap Node<T>*> DoublyLinkedList.find(T value) {
    heap Node<T>* currentNode = this.head;
    while currentNode != nil<heap Node<T>*> {
        // Check condition
        if currentNode.value == value {
            return currentNode;
        }
        // Move to next node
        currentNode = currentNode.next;
    }
    return nil<heap Node<T>*>;
}*/