f<int> main() {
    int[10][10] a;
    for int i = 0; i < row; i++ {
        for int j = 0; j < col; j++ {
            a[i][j] = i * j;
        }
    }
    printf("Cell [1,3]: %d", a[1][3]);
}