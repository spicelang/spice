type Struct struct {
    int _fieldA
    bool _fieldB
    string _fieldC
}

f<int> main() {
    printf("Alignment of double: %d\n", alignof(-19.34989));
    printf("Alignment of int: %d\n", alignof(353));
    printf("Alignment of short: %d\n", alignof(35s));
    printf("Alignment of long: %d\n", alignof(9223372036854775807l));
    printf("Alignment of byte: %d\n", alignof((byte) 13));
    printf("Alignment of char: %d\n", alignof((char) 65));
    printf("Alignment of string: %d\n", alignof("Hello Spice!"));
    printf("Alignment of bool: %d\n", alignof(false));
    printf("Alignment of int[]: %d\n", alignof([1, 2, 3, 4, 5, 6, 7]));
    int intVariable = 123;
    printf("Alignment of int*: %d\n", alignof(&intVariable));
    printf("Alignment of struct instance: %d\n", alignof(type Struct));
}