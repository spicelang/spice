f<int> test(string _input) {
    return 12;
}

f<int> invoke(f<int>(string)** fctPtr) {
    return fctPtr("string");
}

f<int> invoke(f<int>(string)& fctPtr) {
    return fctPtr("string");
}

f<int> main() {
    f<int>(string) testFct = test;
    f<int>(string)* testFctPtr = &testFct;
    printf("%d\n", invoke(&testFctPtr));
    printf("%d\n", invoke(testFct));
}