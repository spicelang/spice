const int MODE_ALL_RWX = 0o0000777;

ext<byte*> malloc(long);
ext free(char*);

f<int> main() {
    byte* address = malloc(1l);
    *address = (byte) 12;
    free(address);
}