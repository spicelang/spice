f<int> main() {
    printf("Hi World!");
}

/*type T int|long;

type TestStruct<T> struct {
    T _f1
    unsigned long length
}

p TestStruct.ctor(const unsigned long initialLength) {
    this.length = initialLength;
}

p TestStruct.printLength() {
    printf("%d\n", this.length);
}

type Alias alias TestStruct<long>;

f<int> main() {
    Alias a = Alias{12345l, (unsigned long) 54321l};
    a.printLength();
    dyn b = Alias(12l);
    b.printLength();
}*/

/*type TestStruct struct {

}

f<int> TestStruct.test(const string& input) {
    printf("%s", input);
    return 1;
}

f<int> test() {
    printf("Hi");
    return 12;
}

f<int> main() {
    TestStruct ts;
    int t = ts.test("Test");
    t = test();
}*/