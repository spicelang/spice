type Visitable interface {
    f<bool> accept<int>(Visitor*);
}

f<int> main() {

}
