f<int> main() {
    assert false;
    /*f<string>() callbackWithoutArgs = () -> string {
        return "Callback called!\n";
    };
    printf("%s", callbackWithoutArgs());

    f<String>(String&, double) callbackWithArgs1 = (String& str, double d) -> String {
        printf("Callback called with args: %s, %f\n", str, d);
        return str;
    };
    printf("%s\n", callbackWithArgs1(String("Hello"), 3.14));

    f<short>(String, short) callbackWithArgs2 = (String str, short b) -> short {
        printf("Callback called with args: %s, %d\n", str, b);
        return ~b;
    };
    printf("%d\n", (callbackWithArgs2(String("Hello World!"), 321s) ^ 956s) == 1 ? 9 : 12);*/
}


/*type T int|long;

type TestStruct<T> struct {
    T _f1
    unsigned long length
}

p TestStruct.ctor(const unsigned long initialLength) {
    this.length = initialLength;
}

p TestStruct.printLength() {
    printf("%d\n", this.length);
}

type Alias alias TestStruct<long>;

f<int> main() {
    Alias a = Alias{12345l, (unsigned long) 54321l};
    a.printLength();
    dyn b = Alias(12l);
    b.printLength();
}*/

/*type TestStruct struct {
    long lng
    String str
    int i
}

p TestStruct.dtor() {}

f<TestStruct> fct(int& ref) {
    TestStruct ts = TestStruct{ 6l, String("test string"), ref };
    return ts;
}

f<int> main() {
    int test = 987654;
    const TestStruct res = fct(test);
    printf("Long: %d\n", res.lng);
    printf("String: %s\n", res.str.getRaw());
    printf("Int: %d\n", res.i);
}*/