// Add generic type definitions
type V1 dyn;
type V2 dyn;

/**
 * A pair in Spice is a commonly used data structure, which saves two values of arbitrary type together in a correlation
 */
public type Pair<V1, V2> struct {
    V1 first
    V2 second
}

public inline p Pair.ctor(V1 first, V2 second) {
    this.first = first;
    this.second = second;
}

public inline f<V1&> Pair.getFirst() {
    return this.first;
}

public inline f<V2&> Pair.getSecond() {
    return this.second;
}

public inline p Pair.setFirst(const V1& first) {
    this.first = first;
}

public inline p Pair.setSecond(const V2& second) {
    this.second = second;
}

public f<bool> operator==<V1, V2>(const Pair<V1, V2>& lhs, const Pair<V1, V2>& rhs) {
    return lhs.first == rhs.first && lhs.second == rhs.second;
}

public f<bool> operator!=<V1, V2>(const Pair<V1, V2>& lhs, const Pair<V1, V2>& rhs) {
    return !(lhs == rhs);
}