// Std imports

// Own imports

// Enums
public type SymbolState enum {
    DECLARED,
    INITIALIZED
}

public type SymbolTableEntry struct {

}

public p SymbolTableEntry.ctor() {

}