// Syscall numbers
public const unsigned short SYSCALL_READ                   = 0us;
public const unsigned short SYSCALL_WRITE                  = 1us;
public const unsigned short SYSCALL_OPEN                   = 2us;
public const unsigned short SYSCALL_CLOSE                  = 3us;
public const unsigned short SYSCALL_STAT                   = 4us;
public const unsigned short SYSCALL_FSTAT                  = 5us;
public const unsigned short SYSCALL_LSTAT                  = 6us;
public const unsigned short SYSCALL_POLL                   = 7us;
public const unsigned short SYSCALL_LSEEK                  = 8us;
public const unsigned short SYSCALL_MMAP                   = 9us;
public const unsigned short SYSCALL_MPROTECT               = 10us;
public const unsigned short SYSCALL_MUNMAP                 = 11us;
public const unsigned short SYSCALL_BRK                    = 12us;
public const unsigned short SYSCALL_RT_SIGACTION           = 13us;
public const unsigned short SYSCALL_RT_SIGPROCMASK         = 14us;
public const unsigned short SYSCALL_RT_SIGRETURN           = 15us;
public const unsigned short SYSCALL_IOCTL                  = 16us;
public const unsigned short SYSCALL_PREAD64                = 17us;
public const unsigned short SYSCALL_PWRITE64               = 18us;
public const unsigned short SYSCALL_READV                  = 19us;
public const unsigned short SYSCALL_WRITEV                 = 20us;
public const unsigned short SYSCALL_ACCESS                 = 21us;
public const unsigned short SYSCALL_PIPE                   = 22us;
public const unsigned short SYSCALL_SELECT                 = 23us;
public const unsigned short SYSCALL_SCHED_YIELD            = 24us;
public const unsigned short SYSCALL_MREMAP                 = 25us;
public const unsigned short SYSCALL_MSYNC                  = 26us;
public const unsigned short SYSCALL_MINCORE                = 27us;
public const unsigned short SYSCALL_MADVISE                = 28us;
public const unsigned short SYSCALL_SHMGET                 = 29us;
public const unsigned short SYSCALL_SHMAT                  = 30us;
public const unsigned short SYSCALL_SHMCTL                 = 31us;
public const unsigned short SYSCALL_DUP                    = 32us;
public const unsigned short SYSCALL_DUP2                   = 33us;
public const unsigned short SYSCALL_PAUSE                  = 34us;
public const unsigned short SYSCALL_NANOSLEEP              = 35us;
public const unsigned short SYSCALL_GETITIMER              = 36us;
public const unsigned short SYSCALL_ALARM                  = 37us;
public const unsigned short SYSCALL_SETITIMER              = 38us;
public const unsigned short SYSCALL_GETPID                 = 39us;
public const unsigned short SYSCALL_SENDFILE               = 40us;
public const unsigned short SYSCALL_SOCKET                 = 41us;
public const unsigned short SYSCALL_CONNECT                = 42us;
public const unsigned short SYSCALL_ACCEPT                 = 43us;
public const unsigned short SYSCALL_SENDTO                 = 44us;
public const unsigned short SYSCALL_RECVFROM               = 45us;
public const unsigned short SYSCALL_SENDMSG                = 46us;
public const unsigned short SYSCALL_RECVMSG                = 47us;
public const unsigned short SYSCALL_SHUTDOWN               = 48us;
public const unsigned short SYSCALL_BIND                   = 49us;
public const unsigned short SYSCALL_LISTEN                 = 50us;
public const unsigned short SYSCALL_GETSOCKNAME            = 51us;
public const unsigned short SYSCALL_GETPEERNAME            = 52us;
public const unsigned short SYSCALL_SOCKETPAIR             = 53us;
public const unsigned short SYSCALL_SETSOCKOPT             = 54us;
public const unsigned short SYSCALL_GETSOCKOPT             = 55us;
public const unsigned short SYSCALL_CLONE                  = 56us;
public const unsigned short SYSCALL_FORK                   = 57us;
public const unsigned short SYSCALL_VFORK                  = 58us;
public const unsigned short SYSCALL_EXECVE                 = 59us;
public const unsigned short SYSCALL_EXIT                   = 60us;
public const unsigned short SYSCALL_WAIT4                  = 61us;
public const unsigned short SYSCALL_KILL                   = 62us;
public const unsigned short SYSCALL_UNAME                  = 63us;
public const unsigned short SYSCALL_SEMGET                 = 64us;
public const unsigned short SYSCALL_SEMOP                  = 65us;
public const unsigned short SYSCALL_SEMCTL                 = 66us;
public const unsigned short SYSCALL_SHMDT                  = 67us;
public const unsigned short SYSCALL_MSGGET                 = 68us;
public const unsigned short SYSCALL_MSGSND                 = 69us;
public const unsigned short SYSCALL_MSGRCV                 = 70us;
public const unsigned short SYSCALL_MSGCTL                 = 71us;
public const unsigned short SYSCALL_FCNTL                  = 72us;
public const unsigned short SYSCALL_FLOCK                  = 73us;
public const unsigned short SYSCALL_FSYNC                  = 74us;
public const unsigned short SYSCALL_FDATASYNC              = 75us;
public const unsigned short SYSCALL_TRUNCATE               = 76us;
public const unsigned short SYSCALL_FTRUNCATE              = 77us;
public const unsigned short SYSCALL_GETDENTS               = 78us;
public const unsigned short SYSCALL_GETCWD                 = 79us;
public const unsigned short SYSCALL_CHDIR                  = 80us;
public const unsigned short SYSCALL_FCHDIR                 = 81us;
public const unsigned short SYSCALL_RENAME                 = 82us;
public const unsigned short SYSCALL_MKDIR                  = 83us;
public const unsigned short SYSCALL_RMDIR                  = 84us;
public const unsigned short SYSCALL_CREAT                  = 85us;
public const unsigned short SYSCALL_LINK                   = 86us;
public const unsigned short SYSCALL_UNLINK                 = 87us;
public const unsigned short SYSCALL_SYMLINK                = 88us;
public const unsigned short SYSCALL_READLINK               = 89us;
public const unsigned short SYSCALL_CHMOD                  = 90us;
public const unsigned short SYSCALL_FCHMOD                 = 91us;
public const unsigned short SYSCALL_CHOWN                  = 92us;
public const unsigned short SYSCALL_FCHOWN                 = 93us;
public const unsigned short SYSCALL_LCHOWN                 = 94us;
public const unsigned short SYSCALL_UMASK                  = 95us;
public const unsigned short SYSCALL_GETTIMEOFDAY           = 96us;
public const unsigned short SYSCALL_GETRLIMIT              = 97us;
public const unsigned short SYSCALL_GETRUSAGE              = 98us;
public const unsigned short SYSCALL_SYSINFO                = 99us;
public const unsigned short SYSCALL_TIMES                  = 100us;
public const unsigned short SYSCALL_PTRACE                 = 101us;
public const unsigned short SYSCALL_GETUID                 = 102us;
public const unsigned short SYSCALL_SYSLOG                 = 103us;
public const unsigned short SYSCALL_GETGID                 = 104us;
public const unsigned short SYSCALL_SETUID                 = 105us;
public const unsigned short SYSCALL_SETGID                 = 106us;
public const unsigned short SYSCALL_GETEUID                = 107us;
public const unsigned short SYSCALL_GETEGID                = 108us;
public const unsigned short SYSCALL_SETPGID                = 109us;
public const unsigned short SYSCALL_GETPPID                = 110us;
public const unsigned short SYSCALL_GETPGRP                = 111us;
public const unsigned short SYSCALL_SETSID                 = 112us;
public const unsigned short SYSCALL_SETREUID               = 113us;
public const unsigned short SYSCALL_SETREGID               = 114us;
public const unsigned short SYSCALL_GETGROUPS              = 115us;
public const unsigned short SYSCALL_SETGROUPS              = 116us;
public const unsigned short SYSCALL_SETRESUID              = 117us;
public const unsigned short SYSCALL_GETRESUID              = 118us;
public const unsigned short SYSCALL_SETRESGID              = 119us;
public const unsigned short SYSCALL_GETRESGID              = 120us;
public const unsigned short SYSCALL_GETPGID                = 121us;
public const unsigned short SYSCALL_SETFSUID               = 122us;
public const unsigned short SYSCALL_SETFSGID               = 123us;
public const unsigned short SYSCALL_GETSID                 = 124us;
public const unsigned short SYSCALL_CAPGET                 = 125us;
public const unsigned short SYSCALL_CAPSET                 = 126us;
public const unsigned short SYSCALL_RT_SIGPENDING          = 127us;
public const unsigned short SYSCALL_RT_SIGTIMEDWAIT        = 128us;
public const unsigned short SYSCALL_RT_SIGQUEUEINFO        = 129us;
public const unsigned short SYSCALL_RT_SIGSUSPEND          = 130us;
public const unsigned short SYSCALL_SIGALTSTACK            = 131us;
public const unsigned short SYSCALL_UTIME                  = 132us;
public const unsigned short SYSCALL_MKNOD                  = 133us;
public const unsigned short SYSCALL_USELIB                 = 134us;
public const unsigned short SYSCALL_PERSONALITY            = 135us;
public const unsigned short SYSCALL_USTAT                  = 136us;
public const unsigned short SYSCALL_STATFS                 = 137us;
public const unsigned short SYSCALL_FSTATFS                = 138us;
public const unsigned short SYSCALL_SYSFS                  = 139us;
public const unsigned short SYSCALL_GETPRIORITY            = 140us;
public const unsigned short SYSCALL_SETPRIORITY            = 141us;
public const unsigned short SYSCALL_SCHED_SETPARAM         = 142us;
public const unsigned short SYSCALL_SCHED_GETPARAM         = 143us;
public const unsigned short SYSCALL_SCHED_SETSCHEDULER     = 144us;
public const unsigned short SYSCALL_SCHED_GETSCHEDULER     = 145us;
public const unsigned short SYSCALL_SCHED_GET_PRIORITY_MAX = 146us;
public const unsigned short SYSCALL_SCHED_GET_PRIORITY_MIN = 147us;
public const unsigned short SYSCALL_SCHED_RR_GET_INTERVAL  = 148us;
public const unsigned short SYSCALL_MLOCK                  = 149us;
public const unsigned short SYSCALL_MUNLOCK                = 150us;
public const unsigned short SYSCALL_MLOCKALL               = 151us;
public const unsigned short SYSCALL_MUNLOCKALL             = 152us;
public const unsigned short SYSCALL_VHANGUP                = 153us;
public const unsigned short SYSCALL_MODIFY_LDT             = 154us;
public const unsigned short SYSCALL_PIVOT_ROOT             = 155us;
public const unsigned short SYSCALL__SYSCTL                = 156us;
public const unsigned short SYSCALL_PRCTL                  = 157us;
public const unsigned short SYSCALL_ARCH_PRCTL             = 158us;
public const unsigned short SYSCALL_ADJTIMEX               = 159us;
public const unsigned short SYSCALL_SETRLIMIT              = 160us;
public const unsigned short SYSCALL_CHROOT                 = 161us;
public const unsigned short SYSCALL_SYNC                   = 162us;
public const unsigned short SYSCALL_ACCT                   = 163us;
public const unsigned short SYSCALL_SETTIMEOFDAY           = 164us;
public const unsigned short SYSCALL_MOUNT                  = 165us;
public const unsigned short SYSCALL_UMOUNT2                = 166us;
public const unsigned short SYSCALL_SWAPON                 = 167us;
public const unsigned short SYSCALL_SWAPOFF                = 168us;
public const unsigned short SYSCALL_REBOOT                 = 169us;
public const unsigned short SYSCALL_SETHOSTNAME            = 170us;
public const unsigned short SYSCALL_SETDOMAINNAME          = 171us;
public const unsigned short SYSCALL_IOPL                   = 172us;
public const unsigned short SYSCALL_IOPERM                 = 173us;
public const unsigned short SYSCALL_CREATE_MODULE          = 174us;
public const unsigned short SYSCALL_INIT_MODULE            = 175us;
public const unsigned short SYSCALL_DELETE_MODULE          = 176us;
public const unsigned short SYSCALL_GET_KERNEL_SYMS        = 177us;
public const unsigned short SYSCALL_QUERY_MODULE           = 178us;
public const unsigned short SYSCALL_QUOTACTL               = 179us;
public const unsigned short SYSCALL_NFSSERVCTL             = 180us;
public const unsigned short SYSCALL_GETPMSG                = 181us;
public const unsigned short SYSCALL_PUTPMSG                = 182us;
public const unsigned short SYSCALL_AFS_SYSCALL            = 183us;
public const unsigned short SYSCALL_TUXCALL                = 184us;
public const unsigned short SYSCALL_SECURITY               = 185us;
public const unsigned short SYSCALL_GETTID                 = 186us;
public const unsigned short SYSCALL_READAHEAD              = 187us;
public const unsigned short SYSCALL_SETXATTR               = 188us;
public const unsigned short SYSCALL_LSETXATTR              = 189us;
public const unsigned short SYSCALL_FSETXATTR              = 190us;
public const unsigned short SYSCALL_GETXATTR               = 191us;
public const unsigned short SYSCALL_LGETXATTR              = 192us;
public const unsigned short SYSCALL_FGETXATTR              = 193us;
public const unsigned short SYSCALL_LISTXATTR              = 194us;
public const unsigned short SYSCALL_LLISTXATTR             = 195us;
public const unsigned short SYSCALL_FLISTXATTR             = 196us;
public const unsigned short SYSCALL_REMOVEXATTR            = 197us;
public const unsigned short SYSCALL_LREMOVEXATTR           = 198us;
public const unsigned short SYSCALL_FREMOVEXATTR           = 199us;
public const unsigned short SYSCALL_TKILL                  = 200us;
public const unsigned short SYSCALL_TIME                   = 201us;
public const unsigned short SYSCALL_FUTEX                  = 202us;
public const unsigned short SYSCALL_SCHED_SETAFFINITY      = 203us;
public const unsigned short SYSCALL_SCHED_GETAFFINITY      = 204us;
public const unsigned short SYSCALL_SET_THREAD_AREA        = 205us;
public const unsigned short SYSCALL_IO_SETUP               = 206us;
public const unsigned short SYSCALL_IO_DESTROY             = 207us;
public const unsigned short SYSCALL_IO_GETEVENTS           = 208us;
public const unsigned short SYSCALL_IO_SUBMIT              = 209us;
public const unsigned short SYSCALL_IO_CANCEL              = 210us;
public const unsigned short SYSCALL_GET_THREAD_AREA        = 211us;
public const unsigned short SYSCALL_LOOKUP_DCOOKIE         = 212us;
public const unsigned short SYSCALL_EPOLL_CREATE           = 213us;
public const unsigned short SYSCALL_EPOLL_CTL_OLD          = 214us;
public const unsigned short SYSCALL_EPOLL_WAIT_OLD         = 215us;
public const unsigned short SYSCALL_REMAP_FILE_PAGES       = 216us;
public const unsigned short SYSCALL_GETDENTS64             = 217us;
public const unsigned short SYSCALL_SET_TID_ADDRESS        = 218us;
public const unsigned short SYSCALL_RESTART_SYSCALL        = 219us;
public const unsigned short SYSCALL_SEMTIMEDOP             = 220us;
public const unsigned short SYSCALL_FADVISE64              = 221us;
public const unsigned short SYSCALL_TIMER_CREATE           = 222us;
public const unsigned short SYSCALL_TIMER_SETTIME          = 223us;
public const unsigned short SYSCALL_TIMER_GETTIME          = 224us;
public const unsigned short SYSCALL_TIMER_GETOVERRUN       = 225us;
public const unsigned short SYSCALL_TIMER_DELETE           = 226us;
public const unsigned short SYSCALL_CLOCK_SETTIME          = 227us;
public const unsigned short SYSCALL_CLOCK_GETTIME          = 228us;
public const unsigned short SYSCALL_CLOCK_GETRES           = 229us;
public const unsigned short SYSCALL_CLOCK_NANOSLEEP        = 230us;
public const unsigned short SYSCALL_EXIT_GROUP             = 231us;
public const unsigned short SYSCALL_EPOLL_WAIT             = 232us;
public const unsigned short SYSCALL_EPOLL_CTL              = 233us;
public const unsigned short SYSCALL_TGKILL                 = 234us;
public const unsigned short SYSCALL_UTIMES                 = 235us;
public const unsigned short SYSCALL_VSERVER                = 236us;
public const unsigned short SYSCALL_MBIND                  = 237us;
public const unsigned short SYSCALL_SET_MEMPOLICY          = 238us;
public const unsigned short SYSCALL_GET_MEMPOLICY          = 239us;
public const unsigned short SYSCALL_MQ_OPEN                = 240us;
public const unsigned short SYSCALL_MQ_UNLINK              = 241us;
public const unsigned short SYSCALL_MQ_TIMEDSEND           = 242us;
public const unsigned short SYSCALL_MQ_TIMEDRECEIVE        = 243us;
public const unsigned short SYSCALL_MQ_NOTIFY              = 244us;
public const unsigned short SYSCALL_MQ_GETSETATTR          = 245us;
public const unsigned short SYSCALL_KEXEC_LOAD             = 246us;
public const unsigned short SYSCALL_WAITID                 = 247us;
public const unsigned short SYSCALL_ADD_KEY                = 248us;
public const unsigned short SYSCALL_REQUEST_KEY            = 249us;
public const unsigned short SYSCALL_KEYCTL                 = 250us;
public const unsigned short SYSCALL_IOPRIO_SET             = 251us;
public const unsigned short SYSCALL_IOPRIO_GET             = 252us;
public const unsigned short SYSCALL_INOTIFY_INIT           = 253us;
public const unsigned short SYSCALL_INOTIFY_ADD_WATCH      = 254us;
public const unsigned short SYSCALL_INOTIFY_RM_WATCH       = 255us;
public const unsigned short SYSCALL_MIGRATE_PAGES          = 256us;
public const unsigned short SYSCALL_OPENAT                 = 257us;
public const unsigned short SYSCALL_MKDIRAT                = 258us;
public const unsigned short SYSCALL_MKNODAT                = 259us;
public const unsigned short SYSCALL_FCHOWNAT               = 260us;
public const unsigned short SYSCALL_FUTIMESAT              = 261us;
public const unsigned short SYSCALL_NEWFSTATAT             = 262us;
public const unsigned short SYSCALL_UNLINKAT               = 263us;
public const unsigned short SYSCALL_RENAMEAT               = 264us;
public const unsigned short SYSCALL_LINKAT                 = 265us;
public const unsigned short SYSCALL_SYMLINKAT              = 266us;
public const unsigned short SYSCALL_READLINKAT             = 267us;
public const unsigned short SYSCALL_FCHMODAT               = 268us;
public const unsigned short SYSCALL_FACCESSAT              = 269us;
public const unsigned short SYSCALL_PSELECT6               = 270us;
public const unsigned short SYSCALL_PPOLL                  = 271us;
public const unsigned short SYSCALL_UNSHARE                = 272us;
public const unsigned short SYSCALL_SET_ROBUST_LIST        = 273us;
public const unsigned short SYSCALL_GET_ROBUST_LIST        = 274us;
public const unsigned short SYSCALL_SPLICE                 = 275us;
public const unsigned short SYSCALL_TEE                    = 276us;
public const unsigned short SYSCALL_SYNC_FILE_RANGE        = 277us;
public const unsigned short SYSCALL_VMSPLICE               = 278us;
public const unsigned short SYSCALL_MOVE_PAGES             = 279us;
public const unsigned short SYSCALL_UTIMENSAT              = 280us;
public const unsigned short SYSCALL_EPOLL_PWAIT            = 281us;
public const unsigned short SYSCALL_SIGNALFD               = 282us;
public const unsigned short SYSCALL_TIMERFD_CREATE         = 283us;
public const unsigned short SYSCALL_EVENTFD                = 284us;
public const unsigned short SYSCALL_FALLOCATE              = 285us;
public const unsigned short SYSCALL_TIMERFD_SETTIME        = 286us;
public const unsigned short SYSCALL_TIMERFD_GETTIME        = 287us;
public const unsigned short SYSCALL_ACCEPT4                = 288us;
public const unsigned short SYSCALL_SIGNALFD4              = 289us;
public const unsigned short SYSCALL_EVENTFD2               = 290us;
public const unsigned short SYSCALL_EPOLL_CREATE1          = 291us;
public const unsigned short SYSCALL_DUP3                   = 292us;
public const unsigned short SYSCALL_PIPE2                  = 293us;
public const unsigned short SYSCALL_INOTIFY_INIT1          = 294us;
public const unsigned short SYSCALL_PREADV                 = 295us;
public const unsigned short SYSCALL_PWRITEV                = 296us;
public const unsigned short SYSCALL_RT_TGSIGQUEUEINFO      = 297us;
public const unsigned short SYSCALL_PERF_EVENT_OPEN        = 298us;
public const unsigned short SYSCALL_RECVMMSG               = 299us;
public const unsigned short SYSCALL_FANOTIFY_INIT          = 300us;
public const unsigned short SYSCALL_FANOTIFY_MARK          = 301us;
public const unsigned short SYSCALL_PRLIMIT64              = 302us;
public const unsigned short SYSCALL_NAME_TO_HANDLE_AT      = 303us;
public const unsigned short SYSCALL_OPEN_BY_HANDLE_AT      = 304us;
public const unsigned short SYSCALL_CLOCK_ADJTIME          = 305us;
public const unsigned short SYSCALL_SYNCFS                 = 306us;
public const unsigned short SYSCALL_SENDMMSG               = 307us;
public const unsigned short SYSCALL_SETNS                  = 308us;
public const unsigned short SYSCALL_GETCPU                 = 309us;
public const unsigned short SYSCALL_PROCESS_VM_READV       = 310us;
public const unsigned short SYSCALL_PROCESS_VM_WRITEV      = 311us;
public const unsigned short SYSCALL_KCMP                   = 312us;
public const unsigned short SYSCALL_FINIT_MODULE           = 313us;
public const unsigned short SYSCALL_SCHED_SETATTR          = 314us;
public const unsigned short SYSCALL_SCHED_GETATTR          = 315us;
public const unsigned short SYSCALL_RENAMEAT2              = 316us;
public const unsigned short SYSCALL_SECCOMP                = 317us;
public const unsigned short SYSCALL_GETRANDOM              = 318us;
public const unsigned short SYSCALL_MEMFD_CREATE           = 319us;
public const unsigned short SYSCALL_KEXEC_FILE_LOAD        = 320us;
public const unsigned short SYSCALL_BPF                    = 321us;
public const unsigned short SYSCALL_EXECVEAT               = 322us;
public const unsigned short SYSCALL_USERFAULTFD            = 323us;
public const unsigned short SYSCALL_MEMBARRIER             = 324us;
public const unsigned short SYSCALL_MLOCK2                 = 325us;
public const unsigned short SYSCALL_COPY_FILE_RANGE        = 326us;
public const unsigned short SYSCALL_PREADV2                = 327us;
public const unsigned short SYSCALL_PWRITEV2               = 328us;
public const unsigned short SYSCALL_PKEY_MPROCECT          = 329us;
public const unsigned short SYSCALL_PKEY_ALLOC             = 330us;
public const unsigned short SYSCALL_PKEY_FREE              = 331us;
public const unsigned short SYSCALL_STATX                  = 332us;
