type Iterable interface {
    p print();
}

type A struct : Iterable {
    int a
}

p A.print() {
    printf("A: %d\n", this.a);
}

f<int> main() {
    Iterable a = A{5};
    a.print();
}