f<int> test(string input) {
    return 12;
}

f<int> invoke(f<int>(string)** fctPtr) {
    return fctPtr("string");
}

f<int> invoke(f<int>(string)& fctPtr) {
    return fctPtr("string");
}

f<int> main() {
    f<int>(string) testFct = test;
    printf("%d\n", invoke(&&testFct));
    printf("%d\n", invoke(testFct));
}