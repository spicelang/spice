/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec.Vector<pair.Pair<int, string>> pairVector = vec.Vector<pair.Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair.Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

f<int> main() {
    printf("Array1:\n");
    short arraySize1 = 4s;
    int[arraySize1] array1 = {1, 2, 3};
    array1[3] = 0;
    foreach dyn item : array1 {
        printf("Item: %d\n", item);
    }

    printf("Array2:\n");
    long arraySize2 = 2l;
    string[arraySize2] array2;
    array2[0] = "Hello";
    array2[1] = "world";
    foreach dyn item : array2 {
        printf("Item: %s\n", item);
    }

    printf("Array3:\n");
    int arraySize3 = 3;
    int[arraySize3] array3 = {1, arraySize3, arraySize3};
    foreach dyn item : array3 {
        printf("Item: %d\n", item);
    }

    printf("Array4:\n");
    int arraySize4 = 3;
    int[arraySize4] array4;
    array4 = {1, arraySize4, arraySize4};
    foreach dyn item : array4 {
        printf("Item: %d\n", item);
    }
}