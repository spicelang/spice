import "std/io/cli-option";
import "std/text/print";
import "std/type/string";
import "std/data/vector";
import "std/os/os";
import "std/io/filepath";
import "std/text/stringstream";

public type CliSubcommand struct {
    String name
    String description
    CliSubcommand* parent
    String versionString
    String footerString
    p() callback
    Vector<String> aliases
    Vector<CliSubcommand> subcommands
    Vector<CliOption<bool>> boolOptions
    Vector<CliOption<string>> stringOptions
    Vector<CliOption<String>> stringObjOptions
    Vector<CliOption<int>> intOptions
    Vector<CliOption<FilePath>> filePathOptions
    bool allowUnknownOptions = false
}

public p CliSubcommand.ctor(CliSubcommand* parent, const String& versionString, const String& name, const String& description = String("")) {
    this.name = name;
    this.description = description;
    this.versionString = versionString;
    this.parent = parent;
}

f<bool> CliSubcommand.nameOrAliasMatches(const String& name, const Vector<String>& aliases, string input) {
    if name == input {
        return true;
    }
    foreach const String& a : aliases {
        if a == input {
            return true;
        }
    }
    return false;
}

public f<int> CliSubcommand.parse(unsigned int argc, string[] argv, int layer = 1) {
    // Check if we have any arguments
    if argc == layer {
        if this.callback != nil<p()> {
            p() rc = this.callback;
            rc();
        } else {
            this.printHelp(argv, layer);
            return EXIT_CODE_SUCCESS;
        }
    }

    for unsigned int argNo = layer; argNo < argc; argNo++ {
        string arg = argv[argNo];

        // Check for subcommands
        foreach const CliSubcommand& subcommand : this.subcommands {
            if this.nameOrAliasMatches(subcommand.getName(), subcommand.aliases, arg) {
                return subcommand.parse(argc, argv, layer + 1);
            }
        }

        // Check all commonly used flags
        if (arg == "-h" || arg == "--help") { // Help
            this.printHelp(argv, layer);
            return EXIT_CODE_SUCCESS;
        }
        if (arg == "-v" || arg == "--version") { // Version
            printf("%s\n", this.versionString);
            return EXIT_CODE_SUCCESS;
        }

        // Check for options
        foreach const CliOption<bool>& boolOption : this.boolOptions {
            if this.nameOrAliasMatches(boolOption.getName(), boolOption.getAliases(), arg) {
                bool value = true;
                boolOption.setTargetValue(value);
                boolOption.callCallback(value);
                continue 2; // Continue with next argument
            }
        }
        foreach const CliOption<string>& stringOption : this.stringOptions {
            if this.nameOrAliasMatches(stringOption.getName(), stringOption.getAliases(), arg) {
                // get the argument value
                arg = argv[++argNo];

                stringOption.setTargetValue(arg);
                stringOption.callCallback(arg);
                continue 2; // Continue with next argument
            }
        }
        foreach const CliOption<String>& stringObjOption : this.stringObjOptions {
            if this.nameOrAliasMatches(stringObjOption.getName(), stringObjOption.getAliases(), arg) {
                // get the argument value
                arg = argv[++argNo];
                String parsedArg = String(arg);

                stringObjOption.setTargetValue(parsedArg);
                stringObjOption.callCallback(parsedArg);
                continue 2; // Continue with next argument
            }
        }
        foreach const CliOption<int>& intOption : this.intOptions {
            if this.nameOrAliasMatches(intOption.getName(), intOption.getAliases(), arg) {
                // get the argument value
                arg = argv[++argNo];
                int parsedArg = toInt(arg);

                intOption.setTargetValue(parsedArg);
                intOption.callCallback(parsedArg);
                continue 2; // Continue with next argument
            }
        }
        foreach const CliOption<FilePath>& filePathOption : this.filePathOptions {
            if this.nameOrAliasMatches(filePathOption.getName(), filePathOption.getAliases(), arg) {
                // get the argument value
                arg = argv[++argNo];
                FilePath parsedArg = FilePath(arg);

                filePathOption.setTargetValue(parsedArg);
                filePathOption.callCallback(parsedArg);
                continue 2; // Continue with next argument
            }
        }

        // We could not match the argument
        if !this.allowUnknownOptions {
            printf("Unknown argument: %s\n", arg);
            return EXIT_CODE_ERROR;
        }
    }

    return EXIT_CODE_SUCCESS; // Parsing was successful, return success exit code
}

public const f<const String&> CliSubcommand.getName() {
    return this.name;
}

public const f<const String&> CliSubcommand.getDescription() {
    return this.description;
}

public p CliSubcommand.setVersion(const String& versionString) {
    this.versionString = versionString;
}

public p CliSubcommand.setFooter(const String& footerString) {
    this.footerString = footerString;
}

public p CliSubcommand.setCallback(p() callback) {
    this.callback = callback;
}

public p CliSubcommand.allowUnknownOptions() {
    this.allowUnknownOptions = true;
    foreach CliSubcommand& subcommand : this.subcommands {
        subcommand.allowUnknownOptions();
    }
}

public p CliSubcommand.addAlias(string subCommand) {
    this.aliases.pushBack(String(subCommand));
}

public p CliSubcommand.addAlias(const String& subCommand) {
    this.aliases.pushBack(subCommand);
}

public f<CliSubcommand&> CliSubcommand.addSubcommand(string name, string description) {
    this.subcommands.pushBack(CliSubcommand(this, this.versionString, String(name), String(description)));
    return this.subcommands.back();
}

public f<CliSubcommand&> CliSubcommand.addSubcommand(const String& name, const String& description) {
    this.subcommands.pushBack(CliSubcommand(this, this.versionString, name, description));
    return this.subcommands.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<string>&> CliSubcommand.addOption(string name, string& targetVariable, string description) {
    this.stringOptions.pushBack(CliOption<string>(String(name), targetVariable, String(description)));
    return this.stringOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<string>&> CliSubcommand.addOption(const String& name, string& targetVariable, const String& description) {
    this.stringOptions.pushBack(CliOption<string>(name, targetVariable, description));
    return this.stringOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<string>&> CliSubcommand.addOption(string name, p(string&) callback, string description) {
    this.stringOptions.pushBack(CliOption<string>(String(name), callback, String(description)));
    return this.stringOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<string>&> CliSubcommand.addOption(const String& name, p(string&) callback, const String& description) {
    this.stringOptions.pushBack(CliOption<string>(name, callback, description));
    return this.stringOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<String>&> CliSubcommand.addOption(string name, String& targetVariable, string description) {
    this.stringObjOptions.pushBack(CliOption<String>(String(name), targetVariable, String(description)));
    return this.stringObjOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<String>&> CliSubcommand.addOption(const String& name, String& targetVariable, const String& description) {
    this.stringObjOptions.pushBack(CliOption<String>(name, targetVariable, description));
    return this.stringObjOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<String>&> CliSubcommand.addOption(string name, p(String&) callback, string description) {
    this.stringObjOptions.pushBack(CliOption<String>(String(name), callback, String(description)));
    return this.stringObjOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<String>&> CliSubcommand.addOption(const String& name, p(String&) callback, const String& description) {
    this.stringObjOptions.pushBack(CliOption<String>(name, callback, description));
    return this.stringObjOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<int>&> CliSubcommand.addOption(string name, int& targetVariable, string description) {
    this.intOptions.pushBack(CliOption<int>(String(name), targetVariable, String(description)));
    return this.intOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<int>&> CliSubcommand.addOption(const String& name, int& targetVariable, const String& description) {
    this.intOptions.pushBack(CliOption<int>(name, targetVariable, description));
    return this.intOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<int>&> CliSubcommand.addOption(string name, p(int&) callback, string description) {
    this.intOptions.pushBack(CliOption<int>(String(name), callback, String(description)));
    return this.intOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<int>&> CliSubcommand.addOption(const String& name, p(int&) callback, const String& description) {
    this.intOptions.pushBack(CliOption<int>(name, callback, description));
    return this.intOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<FilePath>&> CliSubcommand.addOption(string name, FilePath& targetVariable, string description) {
    this.filePathOptions.pushBack(CliOption<FilePath>(String(name), targetVariable, String(description)));
    return this.filePathOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<FilePath>&> CliSubcommand.addOption(const String& name, FilePath& targetVariable, const String& description) {
    this.filePathOptions.pushBack(CliOption<FilePath>(name, targetVariable, description));
    return this.filePathOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<FilePath>&> CliSubcommand.addOption(string name, p(FilePath&) callback, string description) {
    this.filePathOptions.pushBack(CliOption<FilePath>(String(name), callback, String(description)));
    return this.filePathOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<FilePath>&> CliSubcommand.addOption(const String& name, p(FilePath&) callback, const String& description) {
    this.filePathOptions.pushBack(CliOption<FilePath>(name, callback, description));
    return this.filePathOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<bool>&> CliSubcommand.addFlag(string name, bool& targetVariable, string description) {
    this.boolOptions.pushBack(CliOption<bool>(String(name), targetVariable, String(description)));
    return this.boolOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<bool>&> CliSubcommand.addFlag(const String& name, bool& targetVariable, const String& description) {
    this.boolOptions.pushBack(CliOption<bool>(name, targetVariable, description));
    return this.boolOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<bool>&> CliSubcommand.addFlag(string name, p(bool&) callback, string description) {
    this.boolOptions.pushBack(CliOption<bool>(String(name), callback, String(description)));
    return this.boolOptions.back();
}

#[ignoreUnusedReturnValue]
public f<CliOption<bool>&> CliSubcommand.addFlag(const String& name, p(bool&) callback, const String& description) {
    this.boolOptions.pushBack(CliOption<bool>(name, callback, description));
    return this.boolOptions.back();
}

public p CliSubcommand.printHelpItem() {
    // Print name and aliases
    StringStream ss;
    ss << "  " << this.name;
    foreach const String& subcommandAlias : this.aliases {
        ss << ", " << subcommandAlias;
    }
    printFixedWidth(ss.str(), 25, true);
    // Description
    printFixedWidth(this.description, 85, true);
    lineBreak();
}

p CliSubcommand.printHelp(string[] argv, int layer) {
    // Build subcommand string
    String subcommand = String(argv[0]);
    for int i = 1; i < layer; i++ {
        subcommand += " " + argv[i];
    }

    // Print usage
    printf("%s\n\nUsage: %s [options]\n", this.description, subcommand);
    // Print subcommands
    if !this.subcommands.isEmpty() {
        printf("\nSubcommands:\n");
        foreach const CliSubcommand& subCommand : this.subcommands {
            subCommand.printHelpItem();
        }
    }

    // Print options
    printf("\nOptions:\n");
    if this.stringOptions.getSize() + this.stringObjOptions.getSize() + this.intOptions.getSize() + this.filePathOptions.getSize() > 0 {
        foreach const CliOption<string>& option : this.stringOptions {
            option.printHelpItem();
        }
        foreach const CliOption<int>& option : this.intOptions {
            option.printHelpItem();
        }
    }

    // Print flags
    printf("\nFlags:\n");
    foreach const CliOption<bool>& flag : this.boolOptions {
        flag.printHelpItem();
    }

    // Print help and version flags
    bool target;
    const dyn helpFlag = CliOption<bool>(String("--help,-h"), target, String("Print this help message"));
    helpFlag.printHelpItem();
    const dyn versionFlag = CliOption<bool>(String("--version,-v"), target, String("Print the version of the application"));
    versionFlag.printHelpItem();

    // Print footer
    if !this.footerString.isEmpty() {
        printf("\n%s\n", this.footerString);
    }
}