f<int> main() {
    int[4] testIntArray = [1, 2, 3, 4];
    printf("Array length: %d\n", len(testIntArray));
}