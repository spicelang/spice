// Std imports
import "std/data/vector";

// Own imports
import "bootstrap/util/common-util";
import "bootstrap/symboltablebuilder/type-chain";
import "bootstrap/symboltablebuilder/scope";

public type Type struct {
    Vector<TypeChainElement> typeChain
    bool isBaseTypeSigned
}

p Type.ctor(SuperType superType) {
    this.typeChain.pushBack(TypeChainElement(superType));
}

p Type.ctor(SuperType superType, const String& subType) {
    this.typeChain.pushBack(TypeChainElement(superType, subType));
}

p Type.ctor(SuperType superType, const String& subType, unsigned long typeId, const TypeChainElementData& data, const QualTypeList& templateTypes) {
    this.typeChain.pushBack(TypeChainElement(superType, subType, typeId, data, templateTypes));
}

p Type.ctor(TypeChain typeChain) {
    this.typeChain = typeChain.typeChain;
}

/**
 * Get the super type of the current type
 *
 * @return Super type
 */
public f<SuperType> Type.getSuperType() {
    assert !this.typeChain.isEmpty();
    return this.typeChain.back().superType;
}

/**
 * Get the sub type of the current type
 *
 * @return Sub type
 */
public f<const String&> Type.getSubType() {
    assert !this.typeChain.isEmpty();
    assert(isOneOf([SuperType::TY_STRUCT, SuperType::TY_INTERFACE, SuperType::TY_ENUM, SuperType::TY_GENERIC]));
    return this.typeChain.back().subType;
}

/**
 * Get the array size of the current type
 *
 * @return Array size
 */
public f<unsigned int> Type.getArraySize() {
    assert !this.typeChain.isEmpty();
    assert(isOneOf([SuperType::TY_ARRAY]));
    return this.typeChain.back().data.arraySize;
}

/**
 * Get the body scope of the current type
 *
 * @return Body scope
 */
public f<Scope*> Type.getBodyScope() {
    assert !this.typeChain.isEmpty();
    assert(isOneOf([SuperType::TY_STRUCT, SuperType::TY_INTERFACE, SuperType::TY_ENUM, SuperType::TY_GENERIC]));
    return this.typeChain.back().data.bodyScope;
}

/**
 * Get the pointer type of the current type as a new type
 *
 * @param node AST node for error messages
 * @return Pointer type of the current type
 */
public f<const Type*> Type.toPtr(const ASTNode* node) {
    // ToDo
    return nil<const Type*>;
}
