import "std/data/vector";

f<int> main() {
    Vector<int> pairVector = Vector<int>();
    pairVector.reserve(10l);
    /*pairVector.pushBack(4);
    pairVector.pushBack(2);
    pairVector.pushBack(4);
    pairVector.pushBack(3);
    pairVector.pushBack(1);
    printf("Cap: %d\n", pairVector.getCapacity());
    printf("Size: %d\n", pairVector.getSize());
    pairVector.pushBack(2);
    pairVector.pushBack(2);
    pairVector.pushBack(2);
    printf("Cap: %d\n", pairVector.getCapacity());
    printf("Size: %d\n", pairVector.getSize());
    printf("Val: %d\n", pairVector.get(2));*/
    pairVector.dtor();
}