dyn TEST = true;
dyn INVALID;

f<int> main() {
    printf("Bool: %d", TEST);
}