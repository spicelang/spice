/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

type Nested struct {
    string nested1
    bool* nested2
}

type TestStruct struct {
    signed int* field1
    double field2
    Nested* nested
}

f<int> main() {
    int input = 12;
    bool boolean = true;
    Nested nestedInstance = Nested { "Hello World!", &boolean };
    dyn instance = TestStruct { &input, 46.34, &nestedInstance };
    TestStruct instance1 = instance;
    printf("Field1: %d, field2: %f", *instance.nested.nested2, instance1.field2);
    printf("Output: %s, %p", instance1.nested.nested1, instance.field1);
}