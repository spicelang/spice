#[core.compiler.mangledName = "pthread_self"]
ext f<byte*> pthreadSelf();

f<int> main() {}