type Person struct {
    string firstName
    string lastName
    unsigned int age
}

p birthday(Person* person) {
    person.age++;
}

f<int> main() {
    dyn mike = Person { "Mike", "Miller", 32 };
    printf("Person: %s, %s", mike.lastName, mike.firstName);
    printf("Age before birthday: %d", mike.age);
    birthday(&mike);
    printf("Age after birthday: %d", mike.age);
}