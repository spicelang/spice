f<int> test(int i, int j = 12, string t = "Test") {
    printf("Test: %d, %s", j, t);
    return i;
}

f<int> main() {
    test(1);
    test(1, 3);
}