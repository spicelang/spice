// Std imports
import "std/type/byte";
import "std/data/vector";
import "std/data/unordered-map";
import "std/time/timer";
import "std/io/filepath";

// Own imports
import "bootstrap/ast/ast-nodes";
import "bootstrap/global/global-resource-manager-intf";
import "bootstrap/global/cache-manager";
import "bootstrap/global/runtime-module-manager";
import "bootstrap/exception/error-manager";
import "bootstrap/linker/external-linker-interface";
import "bootstrap/reader/code-loc";
import "bootstrap/util/memory";
import "bootstrap/util/block-allocator";
import "bootstrap/bindings/llvm/llvm" as llvm;
import "bootstrap/source-file";
import "bootstrap/driver";

// Constants
public const string MAIN_FILE_NAME = "root";
public const string LTO_FILE_NAME = "lto-module";

/**
 * The GlobalResourceManager is instantiated at startup of the compiler and serves as distribution point for globally used assets.
 * This component owns all SourceFile instances and AST nodes and therefore is the resource root of the compiler.
 * Other components of the compiler can request the required global resources from the GlobalResourceManager.
 */
public type GlobalResourceManager struct : IGlobalResourceManager {
    public llvm::LLVMContext context
    public llvm::IRBuilder builder
    public llvm::Module ltoModule
    public llvm::TargetMachine targetMachine
    public DefaultMemoryManager memoryManager
    public Vector<String> compileTimeStringValues
    public BlockAllocator<ASTNode> astNodeAlloc // Used to allocate all AST nodes
    public UnorderedMap<String, heap SourceFile*> sourceFiles // The GlobalResourceManager owns all source files
    public Vector<ASTNode*> astNodes
    public CliOptions& cliOptions
    public ExternalLinkerInterface linker
    public CacheManager cacheManager
    public RuntimeModuleManager runtimeModuleManager
    public Timer totalTimer
    public ErrorManager errorManager
    public bool abortCompilation = false
    unsigned long nextCustomTypeId = BYTE_MAX_VALUE + 1l // Start at 256 because all primitive types come first
}

public p GlobalResourceManager.ctor(CliOptions& cliOptions) {
    this.cliOptions = cliOptions;
    this.builder = llvm::IRBuilder(this.context);
    this.astNodeAlloc = BlockAllocator<ASTNode>(this.memoryManager);

    // Initialize the required LLVM targets
    if cliOptions.isNativeTarget {
        llvm::initializeNativeTarget();
        llvm::initializeNativeAsmPrinter();
    } else {
        llvm::initializeAllTargets();
        llvm::initializeAllTargetMCs();
        llvm::initializeAllAsmPrinters();
    }

    // Create target machine for LLVM
    String cpuName = String("generic");
    if cliOptions.isNativeTarget & cliOptions.useCPUFeatures {
        // Retrieve native CPU name and the supported CPU features
        cpuName = String(llvm::getHostCPUName());

    }

    // Create lto module
    if cliOptions.useLTO {
        this.ltoModule = llvm::Module(LTO_FILE_NAME, this.context);
    }
}

public p GlobalResourceManager.dtor() {
    // Cleanup all statics
    // ToDo: Implement
    // Cleanup all LLVM statics
    llvm::llvm_shutdown();
}

public f<heap SourceFile*> GlobalResourceManager.createSourceFile(SourceFile* parent, const String& depName, const FilePath& path, bool isStdFile) {
    // Check if the source file was already added (e.g. by another source file that imports it)
    const String filePathStr = String(path.toString());

    // Create the new source file if it does not exist yet
    if !this.sourceFiles.contains(filePathStr) {
        //heap SourceFile* newSourceFile = new SourceFile(*this, parent, depName, path, isStdFile);
        //this.sourceFiles.insert(filePathStr, newSourceFile);
    }

    return this.sourceFiles.get(filePathStr);
}

public f<unsigned long> GlobalResourceManager.getNextCustomTypeId() {
    return this.nextCustomTypeId++;
}

public f<unsigned long> GlobalResourceManager.getTotalLineCount() {
    result = 0l;
    /*foreach const SourceFile* sourceFile : sourceFiles {
        result += sourceFile.value.getLineCount();
    }*/
}