type T int|dyn|double;

f<int> foo<T>(T t) {
    return 1;
}

f<int> main() {
    foo(1);
    foo(1.0);
    foo("test");
}