import "source1" as s1;
import "source2" as s2;

f<int> dummy() {
    return 0;
}

f<int> main() {}