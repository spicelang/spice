type T int|long|short;

type CompareResult enum {
    LESS,
    EQUAL,
    GREATER
}

type Compareable<T> interface {
    f<CompareResult> compare<T>(const T&, const T&);
}

type Person struct : Compareable<long> {
    string firstName
    string lastName
    unsigned int age
}

p Person.ctor(string firstName, string lastName, unsigned int age) {
    this.firstName = firstName;
    this.lastName = lastName;
    this.age = age;
}

f<CompareResult> Person.compare(const long& a, const long& b) {
    if a > b { return CompareResult::GREATER; }
    if a < b { return CompareResult::LESS; }
    return CompareResult::EQUAL;
}

f<int> main() {
    Person mike = Person("Mike", "Miller", 43);
    const bool isEqual = mike.compare(22l, 22l) == CompareResult::EQUAL;
    printf("%d", isEqual);
}

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";

f<int> main() {
    Lexer lexer = Lexer("./file.spice");
    Parser parser = Parser(lexer);
    parser.parse();
}*/