import "std/data/unordered-set";

f<int> main() {
    UnorderedSet<int> set;
    set.insert(1);
    set.insert(2);
    set.insert(3);
    set.insert(2); // Duplicate, should not be added
    assert set.contains(2);
    set.remove(2);
    assert !set.contains(2);
    assert set.contains(1);
    assert set.contains(3);
    assert set.getSize() == 2;
    assert !set.isEmpty();
    set.clear();
    assert set.getSize() == 0;
    assert set.isEmpty();
    printf("All assertions passed!\n");
}