// TEST: --sanitizer=type

f<int> main() {
    long l = 100l;
    unsafe {
       double* ptr = cast<double*>(&l);
       *ptr += 2.0;
    }
}