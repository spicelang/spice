import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    Vector<Pair<int, string>> pairVector = Vector<Pair<int, string>>();
    pairVector.pushBack(Pair<int, string>(0, "Hello"));
    pairVector.pushBack(Pair<int, string>(1, "World"));

    Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!\n", p1.getSecond());
}