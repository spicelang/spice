// TEST: --output-container=lib

f<int> add(int a, int b) {
    return a + b;
}