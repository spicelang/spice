f<int> main() {
    p() callbackWithoutArgs = () -> {
        printf("Callback called!\n");
    };
    callbackWithoutArgs();

    p(String&, double) callbackWithArgs1 = (String& str, double d) -> {
        printf("Callback called with args: %s, %f\n", str, d);
    };
    callbackWithArgs1(String("Hello"), 3.14);

    p(String, bool) callbackWithArgs2 = (String str, bool b) -> {
        printf("Callback called with args: %s, %d\n", str, b);
    };
    callbackWithArgs2(String("Hello World!"), false);
}