// Std imports
import "std/text/stringstream";

// Own imports
import "bootstrap/util/code-loc";

public type LexerErrorType enum {
    TOKENIZING_FAILED
}

/**
 * Custom exception for errors, occurring while parsing
 */
public type ParserError struct {
    string errorMessage
}

/**
 * Constructor: Used in case that the exact code position where the error occurred is known
 *
 * @param codeLoc Code location where the error occurred
 * @param errorType Type of the error
 * @param message Error message suffix
 */
public p ParserError.ctor(const CodeLoc* codeLoc, const LexerErrorType errorType, const string message) {
    StringStream msg;
    msg << "[Error|Lexer] " << codeLoc.toPrettyString() << ": " << this.getMessagePrefix(errorType) << ": " << message;
    this.errorMessage = msg.str();
}

/**
 * Get the prefix of the error message for a particular error
 *
 * @param errorType Type of the error
 * @return Prefix string for the error type
 */
f<string> ParserError.getMessagePrefix(const LexerErrorType errorType) {
    switch errorType {
        case LexerErrorType::TOKENIZING_FAILED: { return "Tokenizing failed"; }
        default: { panic(Error("Unknown error")); }
    }
}