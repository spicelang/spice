import "std/time/delay";
import "std/os/cpu";

/**
 * Mutex for reserving a resource for exclusive access. This is useful for improving thread-safety
 */
public type Mutex struct {
	bool occupied = false
}

/**
 * Acquire the mutex
 */
public p Mutex.acquire() {
	while this.occupied {
		yield();
	}
	this.occupied = true;
}

/**
 * Release the mutex
 */
public p Mutex.release() {
	this.occupied = false;
}

/**
 * LockGuard is a RAII wrapper for Mutex
 */
public type LockGuard struct {
    Mutex& mutex
}

/**
 * Acquire the mutex
 */
public p LockGuard.ctor(Mutex& mutex) {
    this.mutex = mutex;
    this.mutex.acquire();
}

/**
 * Release the mutex
 */
public p LockGuard.dtor() {
    this.mutex.release();
}