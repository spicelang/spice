import "std/type/int" as unused;

f<int> main() {}