// Converts an int to a double
f<double> toDouble(int input) {
    // ToDo: Implement
    return 0.0;
}

// Converts an int to a short
f<short> ToShort(int input) {
    return (short) input;
}

// Converts an int to a long
f<long> ToLong(int input) {
    return (long) input;
}

// Converts an int to a byte
f<byte> ToByte(int input) {
    return (byte) input;
}

// Converts an int to a char
f<char> ToChar(int input) {
    return (char) input;
}

// Converts an int to a string
f<string> toString(int input) {
    // ToDo: Implement (See https://github.com/golang/go/blob/master/src/strconv/itoa.go)
    return "";
}

// Converts an int to a boolean
f<bool> toBool(int input) {
    return input >= 1;
}