p testProc(int[4]*** nums) {
    int[4]* nums1 = **nums;
    int[4] nums2 = *nums1;
    nums2[2] = 10;
    printf("1: %d\n", nums2[0]);
    printf("2: %d\n", nums2[1]);
    printf("3: %d\n", nums2[2]);
    printf("4: %d\n", nums2[3]);
}

f<int> main() {
    int[4] intArray = { 1, 2, 3, 4 };
    printf("1: %d\n", intArray[1]);
    testProc(& & &intArray);
}