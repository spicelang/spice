// Syscall numbers
public const unsigned short SYSCALL_IO_SETUP                = 0us;
public const unsigned short SYSCALL_IO_DESTROY              = 1us;
public const unsigned short SYSCALL_IO_SUBMIT               = 2us;
public const unsigned short SYSCALL_IO_CANCEL               = 3us;
public const unsigned short SYSCALL_IO_GETEVENTS            = 4us;
public const unsigned short SYSCALL_SETXATTR                = 5us;
public const unsigned short SYSCALL_LSETXATTR               = 6us;
public const unsigned short SYSCALL_FSETXATTR               = 7us;
public const unsigned short SYSCALL_GETXATTR                = 8us;
public const unsigned short SYSCALL_LGETXATTR               = 9us;
public const unsigned short SYSCALL_FGETXATTR               = 10us;
public const unsigned short SYSCALL_LISTXATTR               = 11us;
public const unsigned short SYSCALL_LLISTXATTR              = 12us;
public const unsigned short SYSCALL_FLISTXATTR              = 13us;
public const unsigned short SYSCALL_REMOVEXATTR             = 14us;
public const unsigned short SYSCALL_LREMOVEXATTR            = 15us;
public const unsigned short SYSCALL_FREMOVEXATTR            = 16us;
public const unsigned short SYSCALL_GETCWD                  = 17us;
public const unsigned short SYSCALL_LOOKUP_DCOOKIE          = 18us;
public const unsigned short SYSCALL_EVENTFD2                = 19us;
public const unsigned short SYSCALL_EPOLL_CREATE1           = 20us;
public const unsigned short SYSCALL_EPOLL_CTL               = 21us;
public const unsigned short SYSCALL_EPOLL_PWAIT             = 22us;
public const unsigned short SYSCALL_DUP                     = 23us;
public const unsigned short SYSCALL_DUP3                    = 24us;
public const unsigned short SYSCALL_FCNTL                   = 25us;
public const unsigned short SYSCALL_INOTIFY_INIT1           = 26us;
public const unsigned short SYSCALL_INOTIFY_ADD_WATCH       = 27us;
public const unsigned short SYSCALL_INOTIFY_RM_WATCH        = 28us;
public const unsigned short SYSCALL_IOCTL                   = 29us;
public const unsigned short SYSCALL_IOPRIO_SET              = 30us;
public const unsigned short SYSCALL_IOPRIO_GET              = 31us;
public const unsigned short SYSCALL_FLOCK                   = 32us;
public const unsigned short SYSCALL_MKNODAT                 = 33us;
public const unsigned short SYSCALL_MKDIRAT                 = 34us;
public const unsigned short SYSCALL_UNLINKAT                = 35us;
public const unsigned short SYSCALL_SYMLINKAT               = 36us;
public const unsigned short SYSCALL_LINKAT                  = 37us;
public const unsigned short SYSCALL_RENAMEAT                = 38us;
public const unsigned short SYSCALL_UMOUNT2                 = 39us;
public const unsigned short SYSCALL_MOUNT                   = 40us;
public const unsigned short SYSCALL_PIVOT_ROOT              = 41us;
public const unsigned short SYSCALL_NFSSERVCTL              = 42us;
public const unsigned short SYSCALL_STATFS                  = 43us;
public const unsigned short SYSCALL_FSTATFS                 = 44us;
public const unsigned short SYSCALL_TRUNCATE                = 45us;
public const unsigned short SYSCALL_FTRUNCATE               = 46us;
public const unsigned short SYSCALL_FALLOCATE               = 47us;
public const unsigned short SYSCALL_FACCESSAT               = 48us;
public const unsigned short SYSCALL_CHDIR                   = 49us;
public const unsigned short SYSCALL_FCHDIR                  = 50us;
public const unsigned short SYSCALL_CHROOT                  = 51us;
public const unsigned short SYSCALL_FCHMOD                  = 52us;
public const unsigned short SYSCALL_FCHMODAT                = 53us;
public const unsigned short SYSCALL_FCHOWNAT                = 54us;
public const unsigned short SYSCALL_FCHOWN                  = 55us;
public const unsigned short SYSCALL_OPENAT                  = 56us;
public const unsigned short SYSCALL_CLOSE                   = 57us;
public const unsigned short SYSCALL_VHANGUP                 = 58us;
public const unsigned short SYSCALL_PIPE2                   = 59us;
public const unsigned short SYSCALL_QUOTACTL                = 60us;
public const unsigned short SYSCALL_GETDENTS64              = 61us;
public const unsigned short SYSCALL_LSEEK                   = 62us;
public const unsigned short SYSCALL_READ                    = 63us;
public const unsigned short SYSCALL_WRITE                   = 64us;
public const unsigned short SYSCALL_READV                   = 65us;
public const unsigned short SYSCALL_WRITEV                  = 66us;
public const unsigned short SYSCALL_PREAD64                 = 67us;
public const unsigned short SYSCALL_PWRITE64                = 68us;
public const unsigned short SYSCALL_PREADV                  = 69us;
public const unsigned short SYSCALL_PWRITEV                 = 70us;
public const unsigned short SYSCALL_SENDFILE                = 71us;
public const unsigned short SYSCALL_PSELECT6                = 72us;
public const unsigned short SYSCALL_PPOLL                   = 73us;
public const unsigned short SYSCALL_SIGNALFD4               = 74us;
public const unsigned short SYSCALL_VMSPLICE                = 75us;
public const unsigned short SYSCALL_SPLICE                  = 76us;
public const unsigned short SYSCALL_TEE                     = 77us;
public const unsigned short SYSCALL_READLINKAT              = 78us;
public const unsigned short SYSCALL_FSTATAT                 = 79us;
public const unsigned short SYSCALL_FSTAT                   = 80us;
public const unsigned short SYSCALL_SYNC                    = 81us;
public const unsigned short SYSCALL_FSYNC                   = 82us;
public const unsigned short SYSCALL_FDATASYNC               = 83us;
public const unsigned short SYSCALL_SYNC_FILE_RANGE         = 84us;
public const unsigned short SYSCALL_TIMERFD_CREATE          = 85us;
public const unsigned short SYSCALL_TIMERFD_SETTIME         = 86us;
public const unsigned short SYSCALL_TIMERFD_GETTIME         = 87us;
public const unsigned short SYSCALL_UTIMENSAT               = 88us;
public const unsigned short SYSCALL_ACCT                    = 89us;
public const unsigned short SYSCALL_CAPGET                  = 90us;
public const unsigned short SYSCALL_CAPSET                  = 91us;
public const unsigned short SYSCALL_PERSONALITY             = 92us;
public const unsigned short SYSCALL_EXIT                    = 93us;
public const unsigned short SYSCALL_EXIT_GROUP              = 94us;
public const unsigned short SYSCALL_WAITID                  = 95us;
public const unsigned short SYSCALL_SET_TID_ADDRESS         = 96us;
public const unsigned short SYSCALL_UNSHARE                 = 97us;
public const unsigned short SYSCALL_FUTEX                   = 98us;
public const unsigned short SYSCALL_SET_ROBUST_LIST         = 99us;
public const unsigned short SYSCALL_GET_ROBUST_LIST         = 100us;
public const unsigned short SYSCALL_NANOSLEEP               = 101us;
public const unsigned short SYSCALL_GETITIMER               = 102us;
public const unsigned short SYSCALL_SETITIMER               = 103us;

// ToDo: Incomplete
