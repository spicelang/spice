/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/data/vector" as vector;

f<int> main() {
    dyn v = vector.Vector<int>{};
    v.push(4);
    v.push(2);
}*/

/*f<int> testFunc(string param = "Test") {
    printf("Test func %s\n", param);
    return 2;
}

f<int> main() {
    int res = testFunc();
    printf("Result: %d\n", res);
}*/

p testProc(int[]*** nums) {
    /*int[]* nums1 = **nums;
    int[] nums2 = *nums1;
    nums2[2] = 10;
    printf("1: %d\n", nums2[0]);
    printf("2: %d\n", nums2[1]);
    printf("3: %d\n", nums2[2]);
    printf("4: %d\n", nums2[3]);*/
}

f<int> main() {
    int[4] intArray = { 1, 2, 3, 4 };
    printf("1: %d\n", intArray[1]);
    testProc(&&&intArray);
}