import "std/data/vector";

import "bootstrap/util/common-util";
import "bootstrap/source-file-intf";

type MockSourceFile struct : ISourceFile {
    string fileName
    unsigned long lineCount = 0l
}

p MockSourceFile.ctor(string fileName, unsigned long lineCount = 0l) {
    this.fileName = fileName;
    this.lineCount = lineCount;
}

f<unsigned long> MockSourceFile.getLineCount() {
    return this.lineCount;
}

f<string> MockSourceFile.getFileName() {
    return this.fileName;
}

f<bool> MockSourceFile.isStdFile() {
    return false;
}

f<int> main() {
    // getLastFragment
    String lastFragment = getLastFragment(String("this.is.a.test.haystack"), ".");
    printf("%s", lastFragment);
    assert lastFragment == "haystack";
    lastFragment = getLastFragment(String(""), ";");
    assert lastFragment == "";
    lastFragment = getLastFragment(String("x-y-z-"), "-");
    assert lastFragment == "";
    // getCircularImportMessage
    const MockSourceFile msf1 = MockSourceFile("file1.spice", 1l);
    const MockSourceFile msf2 = MockSourceFile("file2.spice", 12l);
    const MockSourceFile msf3 = MockSourceFile("file3.spice", 123l);
    const MockSourceFile msf4 = MockSourceFile("file4.spice", 1234l);
    Vector<const ISourceFile*> sourceFiles;
    unsafe {
        sourceFiles.pushBack((const ISourceFile*) &msf1);
        sourceFiles.pushBack((const ISourceFile*) &msf2);
        sourceFiles.pushBack((const ISourceFile*) &msf3);
        sourceFiles.pushBack((const ISourceFile*) &msf4);
    }
    const String cim = getCircularImportMessage(sourceFiles);
    printf("Circular error message:\n%s\n", cim);
    // buildVersionInfo
    const String versionInfo = buildVersionInfo();
    printf("Version info:\n%s\n", versionInfo);

    printf("All assertions passed!");
}