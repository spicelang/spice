import "std/data/map";

f<int> main() {
    Map<int, string> map;
    assert map.getSize() == 0l;
    assert map.isEmpty();
    map.insert(1, "Hello");
    assert map.getSize() == 1l;
    assert !map.isEmpty();
    map.insert(2, "World");
    assert map.getSize() == 2l;
    map.insert(3, "Foo");
    assert map.getSize() == 3l;
    map.insert(4, "Bar");
    assert map.getSize() == 4l;
    assert map.contains(1);
    assert map.contains(2);
    assert map.contains(3);
    assert map.contains(4);
    assert map.get(1) == "Hello";
    assert map.get(2) == "World";
    assert map.get(3) == "Foo";
    assert map.get(4) == "Bar";
    map.remove(2);
    assert map.getSize() == 3l;
    assert !map.contains(2);
    assert !map.isEmpty();
    map.remove(1);
    assert map.getSize() == 2l;
    assert !map.contains(1);
    assert !map.isEmpty();
    string& foo = map.get(3);
    assert foo == "Foo";
    foo = "Baz";
    assert map.get(3) == "Baz";
    Result<string> bar = map.getSafe(4);
    assert bar.isOk();
    assert bar.unwrap() == "Bar";
    Result<string> baz = map.getSafe(5);
    assert baz.isErr();
    map.remove(3);
    assert map.getSize() == 1l;
    assert !map.contains(3);
    assert !map.isEmpty();
    map.remove(4);
    assert map.getSize() == 0l;
    assert !map.contains(4);
    assert map.isEmpty();
}

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";
import "../../src-bootstrap/ast/ast-nodes";

f<int> main() {
    Lexer lexer = Lexer("./test-file.spice");
    Parser parser = Parser(lexer);
    ASTEntryNode* entryNode = parser.parse();
}*/

/*f<int> main() {
    int i = 123; // Captured by ref
    int j = 321; // Captured by val
    dyn lambda = p() {
        printf("Hello from inside: %d\n", i);
        i++;
        i += j;
        printf("Hello from inside: %d\n", i);
    };
    lambda();
    printf("Hello from outside: %d\n", i);
}*/

/*type Visitable interface {
    p print();
}

type Test1 struct : Visitable {
    int f1
}

p Test1.print() {
    printf("Foo: %d", this.f1);
}

f<int> main() {
    Test1 t1 = Test1{123};
    Visitable* v = &t1;
    v.print();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";

f<int> main() {
    Lexer lexer = Lexer("./file.spice");
    Parser parser = Parser(lexer);
    parser.parse();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "std/time/timer";

f<int> main() {
    Timer timer = Timer();
    timer.start();
    Lexer lexer = Lexer("./file.spice");
    unsigned long i = 1l;
    while (!lexer.isEOF()) {
        Token token = lexer.getToken();
        //printf("Token %d: ", i);
        //token.print();
        lexer.advance();
        i++;
    }
    timer.stop();
    printf("Tokens: %d, Time: %d\n", i, timer.getDurationInMillis());
}*/