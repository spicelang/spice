import "os-test2" as s1;

f<int> dummy() {
    return s1::dummy() + dummy();
}

f<int> main() {
    dummy();
}