// This is a test comment
f<int> testFunction(double doubleParam) {
    /*int number;
    number = 123;
    result = number | 5;

    const int testInt = 0;
    double testDouble = 1.5;

    while testDouble < 2.5 {
        for int i = 12; i < 15; i+=2 {
            result = 12;
        }
        testDouble += 2.0;
    }*/
    return 0;
}

p testProcedure(string stringParam, bool boolParam = false) {
    /* Test
    block
    comment */
    /*string testString = "";
    bool testBool = true;
    double result = testString == "" || testBool ? 5.0 : 1.4;
    if result == 5.0 { result = 3.0; }
    int result1 = testFunction(3.0);*/
}

f<int> main() {
    testProcedure("test", true);
    return 0;
}