type Struct struct {
    int& ref
}

f<int> main() {
    int i = 123;
    Struct str = Struct { i }; // test 123
    str.ref = 1234;
    printf("%d, %d", str.ref, i);
}