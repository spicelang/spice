/*int test1 = 10;
//string test2 = "test string";
double test3 = 5.83;
bool test4 = true;

f<int> main() {
    test1 = 11;
    //test2 = "test";
    test3 = 5.84;
    //test4 = false;
    printf("Variable values: %d, %f, %d", test4, test3, test1);
}*/

import "std/type/convert";
import "test/functions";

f<int> main() {
    printf("Test\n");
}