import "test" as s;

p test() {
    printf("p: %f", s.getDouble());
}