type Rule struct {
    bool condBit1
    bool condBit2
    bool condBit3
    bool resultBit
}

const Rule[8] RULE_SET = {
    Rule { false, false, false, false },
    Rule { false, false, true, true },
    Rule { false, true, false, true },
    Rule { false, true, true, true },
    Rule { true, false, false, false },
    Rule { true, false, true, true },
    Rule { true, true, false, true },
    Rule { true, true, true, false }
};

f<int> main() {

}