f<int> main() {
    int[7] intArray = { 1, 5, 4, 0, 12, 12345, 9 };
    foreach (const int idx = 2, const int item : intArray) {
        printf("Item for index %d, %d\n", idx, item);
        idx++;
    }
}