p testProcedure() {
    printf("Test");
}

f<int> main() {
    testProcedure();
    double calcResult = testFunction(2);
    printf("Calc result: %d", calcResult);
    return 0;
}

f<double> testFunction(int testArg) {
    return 1.1432;
}