import "std/iterator/iterator";
import "std/data/pair";
import "std/type/error";

// Generic type definitions
type N int|long|short;

/**
 * A NumberIterator in Spice can be used to iterate over a range of numbers
 */
public type NumberIterator<N> struct : IIterator<N> {
    N currentNumber
    N lowerBound // Inclusive
    N upperBound // Inclusive
}

public p NumberIterator.ctor(N lowerBound, N upperBound) {
    if lowerBound > upperBound { panic(Error("Upper bound is below lower bound")); }
    this.currentNumber = lowerBound;
    this.lowerBound = lowerBound;
    this.upperBound = upperBound;
}

/**
 * Returns the current number of the number range
 *
 * @return Reference to the current number
 */
public inline f<N&> NumberIterator.get() {
    return this.currentNumber;
}

/**
 * Returns the current index and the current number of the number range
 *
 * @return Pair of current index and a reference to the current number
 */
public inline f<Pair<unsigned long, N&>> NumberIterator.getIdx() {
    unsigned long idx = (unsigned long) this.currentNumber - this.lowerBound;
    return Pair<unsigned long, N&>(idx, this.currentNumber);
}

/**
 * Check if the iterator is valid
 *
 * @return true or false
 */
public inline f<bool> NumberIterator.isValid() {
    return this.currentNumber <= this.upperBound;
}

/**
 * Returns the current number of the number range and moves the cursor to the next item
 */
public inline p NumberIterator.next() {
    if !this.isValid() { panic(Error("Calling next() on invalid iterator")); }
    this.currentNumber++;
}

/**
 * Advances the cursor by one
 *
 * @param it NumberIterator
 */
public inline p operator++<N>(NumberIterator<N>& it) {
    if it.currentNumber > it.upperBound { panic(Error("Iterator out of bounds")); }
    it.currentNumber++;
}

/**
 * Move the cursor back by one
 *
 * @param it NumberIterator
 */
public inline p operator--<N>(NumberIterator<N>& it) {
    if it.currentNumber <= it.lowerBound { panic(Error("Iterator out of bounds")); }
    it.currentNumber--;
}

/**
 * Advances the cursor by the given offset
 *
 * @param it NumberIterator
 * @param offset Offset
 */
public inline p operator+=<N>(NumberIterator<N>& it, N offset) {
    if it.currentNumber + offset > it.upperBound || it.currentNumber + offset < it.lowerBound { panic(Error("Iterator out of bounds")); }
    it.currentNumber += offset;
}

/**
 * Move the cursor back by the given offset
 *
 * @param it NumberIterator
 * @param offset Offset
 */
public inline p operator-=<N>(NumberIterator<N>& it, N offset) {
    if it.currentNumber - offset > it.upperBound || it.currentNumber - offset < it.lowerBound { panic(Error("Iterator out of bounds")); }
    it.currentNumber -= offset;
}

/**
 * Convenience wrapper for creating a simple number iterator
 */
public inline f<NumberIterator<N>> range<N>(N begin, N end) {
    return NumberIterator<N>(begin, end);
}

/**
 * Convenience wrapper for creating a simple number iterator
 */
public inline f<NumberIterator<N>> iterate<N>(N lowerBound, N upperBound) {
    return NumberIterator<N>(lowerBound, upperBound);
}