f<int> test(bool a, string b) {
    return 0;
}

f<int> main() {
    f<string>(bool, string) fct = test;
}