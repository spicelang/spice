import "std/type/result";
import "std/type/error";

// Add generic type definitions
type T dyn;

/**
 * Node of a DoublyLinkedList
 */
type Node<T> struct {
    T value
    heap Node<T>* prev = nil<heap Node<T>*>
    heap Node<T>* next = nil<heap Node<T>*>
}

p Node.ctor(const T& value) {
    this.value = value;
}

/**
 * A doubly linked list is a common, dynamically resizable data structure to store uniform data in order.
 * It is characterized by the pointer for every item, pointing to the next one and the pointer, pointing
 * to the previous one.
 */
public type DoublyLinkedList<T> struct {
    heap Node<T>* head = nil<heap Node<T>*>
    heap Node<T>* tail = nil<heap Node<T>*>
    unsigned long size = 0l
}

public p DoublyLinkedList.pushBack(const T& value) {
    heap Node<T>* newNode = this.createNode(value);
    if this.isEmpty() {
        this.head = this.tail = newNode;
    } else {
        this.head.next = newNode;
        newNode.prev = this.head;
        this.head = newNode;
    }
    this.size++;
}

public p DoublyLinkedList.pushFront(const T& value) {
    heap Node<T>* newNode = this.createNode(value);
    if this.isEmpty() {
        this.head = this.tail = newNode;
    } else {
        newNode.next = this.tail;
        this.tail.prev = newNode;
        this.tail = newNode;
    }
    this.size++;
}

public p DoublyLinkedList.insertAt(unsigned long idx, const T& value) {
    // Abort if the index is out of bounds
    if idx < 0 || idx > this.size { panic(Error("Access index out of bound")); }

    heap Node<T>* newNode = this.createNode(value);
    if idx == 0 {
        this.pushFront(value);
    } else if idx == this.size {
        this.pushBack(value);
    } else {
        heap Node<T>* curr = this.tail;
        for unsigned long i = 0l; i < idx - 1l; i++ {
            curr = curr.next;
        }
        newNode.next = curr.next;
        newNode.prev = curr;
        curr.next.prev = newNode;
        curr.next = newNode;
        this.size++;
    }
}

public p DoublyLinkedList.remove(const T& valueToRemove) {
    heap Node<T>* curr = this.tail;
    while curr != nil<heap Node<T>*> {
        if curr.value == valueToRemove {
            if curr == this.tail {
                this.tail = curr.next;
                this.tail.prev = nil<heap Node<T>*>;
            } else if curr == this.head {
                this.head = curr.prev;
                this.head.next = nil<heap Node<T>*>;
            } else {
                curr.prev.next = curr.next;
                curr.next.prev = curr.prev;
            }
            this.size--;
            break;
        }
        curr = curr.next;
    }
}

public p DoublyLinkedList.removeAt(unsigned long idx) {
    // Abort if the index is out of bounds
    if idx < 0 || idx >= this.size { panic(Error("Access index out of bound")); }

    heap Node<T>* curr = this.tail;
    for unsigned long i = 0l; i < idx; i++ {
        curr = curr.next;
    }
    if curr == this.tail {
        this.tail = curr.next;
        this.tail.prev = nil<heap Node<T>*>;
    } else if curr == this.head {
        this.head = curr.prev;
        this.head.next = nil<heap Node<T>*>;
    } else {
        curr.prev.next = curr.next;
        curr.next.prev = curr.prev;
    }
    this.size--;
}

public p DoublyLinkedList.removeAt(unsigned int idx) {
    this.removeAt((unsigned long) idx);
}

public p DoublyLinkedList.removeFront() {
    this.removeAt(0l);
}

public p DoublyLinkedList.removeBack() {
    this.removeAt(this.size - 1l);
}

public inline f<unsigned long> DoublyLinkedList.getSize() {
    return this.size;
}

public inline f<bool> DoublyLinkedList.isEmpty() {
    return this.size == 0l;
}

public f<T&> DoublyLinkedList.get(unsigned long idx) {
    // Abort if the index is out of bounds
    if idx < 0 || idx >= this.size { panic(Error("Access index out of bound")); }

    heap Node<T>* curr = this.tail;
    for unsigned long i = 0l; i < idx; i++ {
        curr = curr.next;
    }
    return curr.value;
}

public f<T&> DoublyLinkedList.get(unsigned int idx) {
    return this.get((unsigned long) idx);
}

public inline f<T&> DoublyLinkedList.getFront() {
    if this.isEmpty() { panic(Error("Access index out of bounds")); }
    return this.tail.value;
}

public inline f<T&> DoublyLinkedList.getBack() {
    if this.isEmpty() { panic(Error("Access index out of bounds")); }
    return this.head.value;
}

f<heap Node<T>*> DoublyLinkedList.createNode(const T& value) {
    heap Node<T>* newNode;
    unsafe {
        Result<heap byte*> allocResult = sAlloc(sizeof(type Node<T>));
        newNode = (heap Node<T>*) allocResult.unwrap();
    }
    newNode.value = value;
    newNode.prev = nil<heap Node<T>*>;
    newNode.next = nil<heap Node<T>*>;
    return newNode;
}