ext f<int> usleep(int);

/**
 * Suspends the execution for the given number of milliseconds
 */
public inline p delay(int millis) {
    usleep(millis * 1000);
}