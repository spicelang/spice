import "os" as os;

f<int> main() {
    printf("Os: %s", getOsName());
}