import "std/type/type-conversion";

f<int> main() {
    // toDouble()
    double asDouble1 = toDouble(true);
    assert asDouble1 == 1.0;
    double asDouble2 = toDouble(false);
    assert asDouble2 == 0.0;

    // toInt()
    int asInt1 = toInt(true);
    assert asInt1 == 1;
    int asInt2 = toInt(false);
    assert asInt2 == 0;

    // toShort()
    short asShort1 = toShort(true);
    assert asShort1 == 1s;
    short asShort2 = toShort(false);
    assert asShort2 == 0s;

    // toLong()
    long asLong1 = toLong(true);
    assert asLong1 == 1l;
    long asLong2 = toLong(false);
    assert asLong2 == 0l;

    // toByte()
    byte asByte1 = toByte(true);
    assert asByte1 == cast<byte>(1);
    byte asByte2 = toByte(false);
    assert asByte2 == cast<byte>(0);

    // toString()
    string asString1 = toString(true);
    assert asString1 == "true";
    string asString2 = toString(false);
    assert asString2 == "false";

    printf("All assertions succeeded");
}