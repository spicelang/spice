import "std/type/result";

// Constants
const unsigned long INITIAL_ALLOC_COUNT = 5l;
const unsigned int RESIZE_FACTOR = 2;

/**
 * Heap-allocated builtin String type to enable dynamic modification in contrast
 * to the primitive string type.
 */
public type String struct {
    heap char* contents    // Pointer to the first char
    unsigned long capacity // Allocated number of chars (without null terminator)
    unsigned long length   // Used number of chars
}

// Generic type definitions
type IntLong      int|long;
type IntLongShort int|long|short;
type StrTy        String|string;
type RawStrChar   string|char;
type StrTyChar    String|string|char;

public p String.ctor(const string value = "") {
    this.length = getRawLength(value);
    this.capacity = this.length > INITIAL_ALLOC_COUNT ? this.length * RESIZE_FACTOR : INITIAL_ALLOC_COUNT;

    // Allocate space for the initial number of elements
    unsafe {
        unsigned long requiredBytes = this.capacity + 1l; // +1 because of null terminator
        Result<heap byte*> allocResult = sAlloc(requiredBytes);
        this.contents = (heap char*) allocResult.unwrap();
    }

    // Save initial value
    unsafe {
        for unsigned long i = 0l; i < this.length + 1l; i++ { // +1 because of null terminator
            this.contents[i] = value[i];
        }
    }
}

public p String.ctor(const char value) {
    this.length = 1l;
    this.capacity = INITIAL_ALLOC_COUNT;

    // Allocate space for the initial number of elements
    unsafe {
        unsigned long requiredBytes = this.capacity + 1l; // +1 because of null terminator
        Result<heap byte*> allocResult = sAlloc(requiredBytes);
        this.contents = (heap char*) allocResult.unwrap();
    }

    // Save initial value
    unsafe {
        this.contents[0] = value;
        this.contents[1] = '\0';
    }
}

public p String.ctor(const String& value) {
    this.length = value.length;
    this.capacity = value.capacity;

    // Allocate space
    unsafe {
        unsigned long requiredBytes = this.capacity + 1l; // +1 because of null terminator
        Result<heap byte*> allocResult = sAlloc(requiredBytes);
        this.contents = (heap char*) allocResult.unwrap();
    }

    // Copy the contents from the other string
    unsafe {
        sCopy((heap byte*) value.contents, (heap byte*) this.contents, value.length + 1l); // +1 because of null terminator
    }
}

/**
 * Appends the given string to the current one
 *
 * @param appendix String to be appended
 */
public p String.append(const string appendix) {
    const unsigned long appendixLength = getRawLength(appendix);
    // Check if we need to re-allocate memory
    while this.capacity < this.length + appendixLength {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Save data
    unsafe {
        for unsigned long i = 0l; i < appendixLength + 1l; i++ { // +1 because of null terminator
            this.contents[this.length++] = appendix[i];
        }
    }
    this.length--; // Remove null terminator
}

/**
 * Appends the given String to the current one
 *
 * @param appendix String to be appended
 */
public p String.append(const String& appendix) {
    this.append(appendix.getRaw());
}

/**
 * Appends the given char to the string and resize it if needed
 *
 * @param c Char to append
 */
public p String.append(const char c) {
    // Check if we need to re-allocate memory
    if this.capacity < this.length + 1l {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Insert the char at the right position
    unsafe {
        this.contents[this.length++] = c;
        this.contents[this.length] = '\0';
    }
}

/**
 * Concatenates two strings and returns the result
 *
 * @parem a String a
 * @param b String b
 * @return Concatenated string
 */
public f<String> operator+<StrTy, StrTyChar>(const StrTy& a, const StrTyChar& b) {
    result = String(a);
    result.append(b);
}

/**
 * Concatenates b to the end of a
 *
 * @param a String a
 * @param b String/string/char b
 */
public p operator+=<StrTyChar>(String& a, const StrTyChar& b) {
    a.append(b);
}

/**
 * Concatenates the given string with itself n times.
 *
 * @param str Input string
 * @param n Multiplication operand
 * @return Result string
 */
public f<String> operator*<IntLongShort>(const String& str, const IntLongShort n) {
    // Shortcuts
    if n < 1 { return String(); }
    if n == 1 { return str; }

    // Copy the input string
    result = String(str);
    const unsigned long newLength = n * str.length;
    result.reserve(newLength);

    // Save the value
    unsafe {
        for unsigned long i = 0l; i < newLength; i++ {
            result.contents[i] = str.contents[i % str.length];
        }
        result.contents[newLength] = '\0';
    }
    result.length = newLength;
}

/**
 * Concatenates the given string with itself n times
 *
 * @param n Multiplication operand
 * @param str Input string
 * @return Result string
 */
public f<String> operator*<IntLongShort>(const IntLongShort n, const String& str) {
    return str * n;
}

/**
 * Concatenates this string with itself n times
 *
 * @param str Input string
 * @param n Multiplication operand
 */
public p operator*=<IntLongShort>(String& str, const IntLongShort n) {
    // Cancel if operand is less than 2
    if n < 2 { return; }

    // Reserve new length
    unsigned long newLength = n * str.length;
    str.reserve(newLength);

    // Save the value
    unsafe {
        for unsigned long i = 0l; i < newLength; i++ {
            str.contents[i] = str.contents[i % str.length];
        }
        str.contents[newLength] = '\0';
    }
    str.length = newLength;
}

/**
 * Checks if two strings have the same value
 *
 * @param a First input string
 * @param b Second input string
 * @return Equal or not
 */
public f<bool> operator==(const String& a, const String& b) {
    // Compare sizes
    if a.length != b.length { return false; }

    // Compare contents
    unsafe {
        for unsigned long i = 0l; i < a.length; i++ {
            if a.contents[i] != b.contents[i] {
                return false;
            }
        }
    }

    return true;
}

/**
 * Checks if two strings have not the same value
 *
 * @param a First input string
 * @param b Second input string
 * @return Not equal or not
 */
public f<bool> operator!=(const String& a, const String& b) {
    return !(a == b);
}

/**
 * Get the raw and immutable string from this container instance
 *
 * @return Raw immutable string
 */
public inline f<string> String.getRaw() {
    unsafe {
        return (string) this.contents;
    }
}

/**
 * Retrieve the current length of the string
 *
 * @return Current length of the string
 */
public inline f<long> String.getLength() {
    return this.length;
}

/**
 * Check if the string is empty
 */
public inline f<bool> String.isEmpty() {
    return this.length == 0;
}

/**
 * Retrieve the current capacity of the string
 *
 * @return Current capacity of the string
 */
 public inline f<long> String.getCapacity() {
     return this.capacity;
 }

/**
 * Checks if the string exhausts its capacity
 *
 * @return Full or not full
 */
public inline f<bool> String.isFull() {
    return this.length == this.capacity;
}

/**
 * Replaces the current contents of the string with an empty string
 */
public p String.clear() {
    this.length = 0l;
    unsafe {
        this.contents[0] = '\0';
    }
}

/**
 * Searches for a substring in a string. Returns -1 if the string was not found.
 *
 * @param startIndex Index where to start the search
 * @return Index, where the substring was found / -1
 */
public f<unsigned long> String.find(string needle, unsigned long startIndex = 0l) {
    // Return -1 if the startIndex is out of bounds
    if startIndex >= this.length { return (unsigned long) -1l; }

    const unsigned long needleLength = getRawLength(needle);
    // Return false if the needle is longer than the haystack
    if this.length < needleLength { return (unsigned long) -1l; }

    // Search needle in haystack
    for unsigned long idx = startIndex; idx <= this.length - needleLength; idx++ {
        // Start matching at startIdx
        for unsigned long charIdx = 0l; charIdx < needleLength; charIdx++ {
            unsafe {
                if this.contents[idx + charIdx] != needle[charIdx] {
                    continue 2;
                }
            }
        }
        // Whole string was matched
        return idx;
    }
    return (unsigned long) -1l;
}

/**
 * Searches for a substring in a string. Returns -1 if the string was not found.
 *
 * @param startIndex Index where to start the search
 * @return Index, where the substring was found / -1
 */
public f<unsigned long> String.find(string needle, unsigned int startIndex) {
    return this.find(needle, (unsigned long) startIndex);
}

/**
 * Searches for a substring in a string from the back. Returns -1 if the string was not found.
 *
 * @param startIndex Index where to start the search
 * @return Index, where the substring was found / -1
 */
public f<unsigned long> String.rfind(string needle, unsigned long startIndex = 0l) {
    // Return -1 if the startIndex is out of bounds
    if startIndex >= this.length { return (unsigned long) -1l; }

    const unsigned long needleLength = getRawLength(needle);
    // Return false if the needle is longer than the haystack
    if this.length < needleLength { return (unsigned long) -1l; }

    if startIndex == 0l { startIndex = this.length - needleLength; }

    // Search needle in haystack
    for unsigned long idx = startIndex; idx >= 0; idx-- {
        // Start matching at startIdx
        for unsigned long charIdx = 0l; charIdx < needleLength; charIdx++ {
            unsafe {
                if this.contents[idx + charIdx] != needle[charIdx] {
                    continue 2;
                }
            }
        }
        // Whole string was matched
        return idx;
    }
    return (unsigned long) -1l;
}

/**
 * Searches for a substring in a string from the back. Returns -1 if the string was not found.
 *
 * @param startIndex Index where to start the search
 * @return Index, where the substring was found / -1
 */
public f<unsigned long> String.rfind(string needle, unsigned int startIndex) {
    return this.rfind(needle, (unsigned long) startIndex);
}

/**
 * Checks if the string contains a substring
 *
 * @param needle Substring to search for
 * @return Found or not
 */
public inline f<bool> String.contains(string needle) {
    return this.find(needle) != -1l;
}

/**
 * Reverse the string
 */
public p String.reverse() {
    unsafe {
        for unsigned long i = 0l; i < this.length / 2l; i++ {
            unsigned long currentUpperIdx = this.length - i - 1l;
            this.contents[i] ^= this.contents[currentUpperIdx];
            this.contents[currentUpperIdx] ^= this.contents[i];
            this.contents[i] ^= this.contents[currentUpperIdx];
        }
    }
}

/**
 * Replace occurrence of substring with the replacement string
 *
 * @param needle Substring to replace
 * @param replacement Replacement for the substring
 */
public f<bool> String.replace(
    string needle,
    string replacement,
    unsigned long startIdx = 0l
) {
    // Abort, if needle or replacement are nullptrs
    if (char*) needle == nil<char*> || (char*) replacement == nil<char*> {
        return false;
    }

    // Find occurrence
    startIdx = this.find(needle, startIdx);
    // Return if not found
    if startIdx == -1l { return false; }

    // Calculate metrics
    const unsigned long needleLength = getRawLength(needle);
    const unsigned long replacementLength = getRawLength(replacement);
    const unsigned long suffixLength = this.length - startIdx - needleLength;
    const unsigned long finalLength = this.length - needleLength + replacementLength;

    // Resize the string if required
    while this.capacity < finalLength {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    unsafe {
        // Move the suffix to the left or right
        const heap char* stringAddr = this.contents;
        const heap char* startAddr = stringAddr + startIdx;
        if needleLength != replacementLength {
            const heap char* oldSuffixAddr = startAddr + needleLength;
            const heap char* newSuffixAddr = startAddr + replacementLength;
            sCopy((heap byte*) oldSuffixAddr, (heap byte*) newSuffixAddr, suffixLength + 1); // +1 because of null terminator
        }

        // Replace needle with replacement
        sCopy((heap byte*) replacement, (heap byte*) startAddr, replacementLength);
    }

    // Update length
    this.length = finalLength;

    return true;
}

/**
 * Replace all occurrences of substring with the replacement string
 *
 * @param needle Substring to replace
 * @param replacement Replacement for the substring
 */
public f<unsigned long> String.replaceAll(string needle, string replacement) {
    unsigned long startIdx = 0l;
    unsigned long foundOccurrences = 0l;
    const unsigned long needleLength = getRawLength(needle);
    const unsigned long replacementLength = getRawLength(replacement);

    while startIdx <= this.length - needleLength {
        if !this.replace(needle, replacement, startIdx) {
            break;
        }
        startIdx += replacementLength;
        foundOccurrences++;
    }

    return foundOccurrences;
}

/**
 * Returns the substring of the current string, starting at position `startIndex` with
 * the length of `length`.
 *
 * @param startIndex Substring start index
 * @param length Length of substring
 * @return Substring
 */
public f<String> String.getSubstring<IntLongShort>(unsigned IntLongShort startIdx, long length = -1l) {
    // Return empty string if the length is 0 or the startIndex is out of bounds
    if length == 0l || startIdx >= this.length {
        return String("");
    }

    // Get everything after startIndex if length is -1
    if length == -1l {
        length = this.length - startIdx;
    }

    // Do not exceed original string length
    if startIdx + length > this.length {
        length = this.length - startIdx;
    }

    // Get substring
    String substring = String("");
    substring.reserve(length);
    const unsigned long endIdx = startIdx + length;
    for unsigned long charIndex = (unsigned long) startIdx; charIndex < endIdx; charIndex++ {
        unsafe {
            substring.contents[charIndex - startIdx] = this.contents[charIndex];
        }
    }

    // Terminate string
    unsafe {
        substring.contents[length] = '\0';
    }

    // Return the substring
    return substring;
}

/**
 * Reserves `charCount` items
 *
 * @param charCount Number of chars to reserve for the string
 */
public p String.reserve<IntLongShort>(unsigned IntLongShort charCount) {
    if charCount > this.capacity {
        this.resize(charCount);
    }
}

/**
 * Re-allocates heap space for the string contents
 *
 * @param newLength new length of the string after resizing
 */
p String.resize<IntLongShort>(unsigned IntLongShort newLength) {
    // Allocate the new memory
    unsafe {
        heap char* oldAddress = this.contents;
        unsigned long requiredBytes = newLength + 1; // +1 because of null terminator
        Result<heap byte*> allocResult = sRealloc((heap byte*) oldAddress, requiredBytes);
        this.contents = (heap char*) allocResult.unwrap();
    }
    // Set new capacity
    this.capacity = newLength;
}

// ======================================================= Static functions ======================================================

/**
 * Returns the length of a string
 *
 * @param input Input string
 * @return Length of the input string
 */
public f<unsigned long> getRawLength(string input) {
    result = 0l;
    while input[result] != '\0' {
        result++;
    }
}

/**
 * Checks the equality of two raw strings
 *
 * @param lhs First input raw string
 * @param rhs Second input raw string
 * @return Equality of lhs and rhs
 */
public f<bool> isRawEqual(string lhs, string rhs) {
    unsigned long lhsLength = getRawLength(lhs);
    unsigned long rhsLength = getRawLength(rhs);
    // Return false immediately if length does not match
    if lhsLength != rhsLength { return false; }
    // Compare chars
    for unsigned long i = 0l; i < lhsLength; i++ {
        if lhs[i] != rhs[i] {
            return false;
        }
    }
    return true;
}