// TEST: --target=aarch64-unknown-linux-gnu

import "std/data/vector";
import "std/text/print";

f<int> main() {
    Vector<String> stringVec;
    stringVec.pushBack(String("Hello "));
    stringVec.pushBack(String("World!"));
    foreach String& str : stringVec {
        print(str);
    }
}