import "std/type/type-conversion";

f<int> main() {
    // toInt()
    int asInt = toInt(123.54);
    assert asInt == 123;

    // toShort()
    short asShort = toShort(12.345);
    assert asShort == 12;

    // toLong()
    long asLong = toLong(534569.2345);
    assert asLong == 534569l;

    // toString()
    //String asString = toString(3.14);
    //assert asString.getRaw() == "3.14";

    // toBool()
    bool asBool1 = toBool(1.0);
    assert asBool1 == true;
    bool asBool2 = toBool(0.0);
    assert asBool2 == false;

    printf("All assertions succeeded");
}