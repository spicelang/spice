f<int> main() {
    const int i = 123;
    i = 1234;
    i++;
    i--;
    ++i;
    --i;
    i += 2;
    i -= 2;
    i *= 2;
    i /= 2;
    i %= 2;
    i ^= 3;
    i <<= 2;
    i >>= 2;
}