import "std/iterator/array-iterator";
import "std/iterator/vector-iterator";

// Generic type definitions
type I dyn; // Item type

/**
 * Convenience wrapper for creating a simple array iterator
 */
public inline f<ArrayIterator<I>> array<I>(I* array, unsigned long size) {
    return ArrayIterator<I>(array, size);
}

/**
 * Convenience wrapper for creating a simple vector iterator
 */
public inline f<VectorIterator<I>> iterate<I>(Vector<I>& container) {
    return VectorIterator<I>(container);
}