// Add generic type definitions
type V1 dyn;
type V2 dyn;
type V3 dyn;

/**
 * A triple in Spice is a commonly used data structure, which saves three values of arbitrary type together in a correlation
 */
public type Triple<V1, V2, V3> struct {
    V1 first
    V2 second
    V3 third
}

public inline p Triple.ctor(V1& first, V2& second, V3& third) {
    this.first = first;
    this.second = second;
    this.third = third;
}

public inline f<V1&> Triple.getFirst() {
    return this.first;
}

public inline f<V2&> Triple.getSecond() {
    return this.second;
}

public inline f<V3&> Triple.getThird() {
    return this.third;
}

public inline p Triple.setFirst(V1& first) {
    this.first = first;
}

public inline p Triple.setSecond(V2& second) {
    this.second = second;
}

public inline p Triple.setThird(V3& third) {
    this.third = third;
}

public f<bool> operator==<V1, V2, V3>(const Triple<V1, V2, V3>& lhs, const Triple<V1, V2, V3>& rhs) {
    return lhs.first == rhs.first && lhs.second == rhs.second && lhs.third == rhs.third;
}

public f<bool> operator!=<V1, V2, V3>(const Triple<V1, V2, V3>& lhs, const Triple<V1, V2, V3>& rhs) {
    return !(lhs == rhs);
}