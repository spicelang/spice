f<int> testFunc() {
    return 12345;
}