type TestStruct struct {
    int a
}

p TestStruct.unusedProcedure() {
    printf("Hello World: %d", this.a);
}

f<string> TestStruct.unusedFunction() {
    printf("%d", this.a);
    return "Hello World";
}

f<int> main() {
    TestStruct _ts;
}