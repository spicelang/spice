// Converts a bool to a double
f<double> toDouble(bool input) {
    return input ? 1.0 : 0.0;
}

// Converts a bool to an int
f<int> toInt(bool input) {
    return input ? 1 : 0;
}

// Converts a bool to a byte
f<byte> toByte(bool input) {
    result = input ? 1 : 0;
}

// Converts a bool to a string
f<string> toString(bool input) {
    return input ? "true" : "false";
}