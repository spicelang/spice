type ITest interface {
    p test();
}

type Test struct : ITest {}

p Test.ctor() {}

p Test.test() {
    printf("Test");
}

p testFct(ITest& test) {
    test.test();
}

f<int> main() {
    Test test = Test();
    ITest& itest = test;
    testFct(itest);
    return 0;
}

/*import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

f<int> main() {
    DefaultMemoryManager defaultMemoryManager;
    IMemoryManager* memoryManager = &defaultMemoryManager;
    BlockAllocator<int> allocator = BlockAllocator<int>(memoryManager, 10);
}*/