ext f<heap byte*> malloc(long);
ext p free(heap byte*);

f<int> main() {
    heap byte* address = malloc(1l);
    *address = (byte) 12;
    free(address);
}