f<int> main(int argc, string[] argv) {
    printf("Argc: %d", argc);
    printf("Argv no. 0: %s", argv[0]);
    if (argc > 1) {
        printf("Argv no. 1: %s", argv[1]);
    }
}