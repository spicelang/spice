f<int> main() {
    int i = 0;
    do {
        i += 1;
        printf("i is now at: %d\n", i);
    } while (i < 10);
}