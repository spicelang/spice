import "std/iterators/ranges";

f<int> main() {
    foreach double item : range(1, 5) {
        printf("Item: %f", item);
    }
}