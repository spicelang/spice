f<int> main() {
    p(int, bool) x = p(int x, bool y = false) {
        x++;
    };
    x(1, true);
}