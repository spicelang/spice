import "../../src-bootstrap/lexer/token";
import "../../src-bootstrap/lexer/lexer";

f<int> main() {
    Lexer lexer = Lexer("./test-file.txt");
    Token token = lexer.getToken();
    assert token.tokenType == TokenType::IDENTIFIER;
}

/*import "std/io/file";

f<int> main() {
    // Write file
    Result<File> fileResult = openFile("./test-file.txt", MODE_WRITE);
    assert fileResult.isOk();
    File file = fileResult.unwrap();
    file.write("Hello, world!\n");
    file.close();

    // Read file
    fileResult = openFile("./test-file.txt", MODE_READ);
    assert fileResult.isOk();
    file = fileResult.unwrap();
    String line = file.readLine();
    printf("%s", line);
    assert line.getRaw() == "Hello, world!\n";
    file.close();

    // Append file
    fileResult = openFile("./test-file.txt", MODE_APPEND);
    assert fileResult.isOk();
    file = fileResult.unwrap();
    file.write("Hello, again!\n");
    file.close();

    // Read file
    fileResult = openFile("./test-file.txt", MODE_READ);
    assert fileResult.isOk();
    file = fileResult.unwrap();
    assert file.readLine() == String("Hello, world!\n");
    assert file.readLine() == String("Hello, again!\n");
    file.close();
}*/