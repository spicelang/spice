f<int> testFunc(int input) {
    if (input > 1) {
        printf("true");
        return;
    }
    printf("false");
    return 0;
}

f<int> main() {
    printf("Result: %d", testFunc(1));
}