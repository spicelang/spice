public f<double> abs(double input) {
    return input < 0 ? -input : input;
}

public f<int> abs(int input) {
    return input < 0 ? -input : input;
}

public f<short> abs(short input) {
    return input < 0 ? -input : input;
}

public f<long> abs(long input) {
    return input < 0 ? -input : input;
}