import "std/data/hash-table";

f<int> main() {
    HashTable<int, int> ht;
    ht.insert(1, 2);
    ht.insert(2, 3);
    ht.insert(3, 4);
    ht.insert(4, 5);
    ht.insert(5, 6);
}