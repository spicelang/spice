f<int> main() {
    int test = 12345678901234567890;
}