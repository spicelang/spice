f<int> main() {
    String test;
    test += "Test";
    printf("%s", test);
}