f<int> main() {
    int i = 1;
    int i = 2;
}