import "std/iterator/array-iterator";

f<int> main() {
    int[7] intArray = [ 1, 5, 4, 0, 12, 12345, 9 ];
    foreach const int item : iterate(intArray, len(intArray)) {
        printf("Item: %d\n", item);
    }
}