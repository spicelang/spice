// Inspired by: https://youtu.be/hmMtQe_mYr0

f<int> main() {
    unsigned long dx = 0x357620655410l;
    while dx > 0 {
        printf("%c", cast<char>(0x726F6C6564574820l >> (((dx >>= 4) & 0xFl) << 3)));
    }
}