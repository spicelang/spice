import "std/data/unordered-map";
import "std/data/vector";
import "std/data/pair";
import "std/math/hash";
import "std/text/stringstream";
import "std/type/type-conversion";

// Generic types
type T dyn;

public type Vertex<T> struct : IHashable {
    T value
}

public p Vertex.ctor(const T& value) {
    this.value = value;
}

public f<T&> Vertex.getValue() {
    return this.value;
}

public f<bool> operator==<T>(const Vertex<T>& v1, const Vertex<T>& v2) {
    return v1.value == v2.value;
}

public f<Hash> Vertex.hash() {
    return hash(this.value);
}

/**
 * Graph data structure
 *
 * ToDo: Add time complexities for common operations
 */
public type Graph<T> struct {
    Vector<Vertex<T>> vertices
    UnorderedMap<Vertex<T>, Vector<Vertex<T>*>> adjList
    bool directed
}

public p Graph.ctor(bool directed = true) {
    this.directed = directed;
}

public f<Vertex<T>&> Graph.addVertex(const T& value) {
    this.vertices.pushBack(Vertex<T>(value));
    Vertex<T>& vertex = this.vertices.back();
    this.adjList.upsert(vertex, Vector<Vertex<T>*>());
    return vertex;
}

public p Graph.addEdge(const Vertex<T>& from, const Vertex<T>& to) {
    if !this.adjList.contains(from) || !this.adjList.contains(to) {
        panic(Error("Graph must already contain both given vertices"));
    }

    Vector<Vertex<T>*>& adjListFrom = this.adjList.get(from);
    adjListFrom.pushBack(&to);
    if !this.directed {
        Vector<Vertex<T>*>& adjListTo = this.adjList.get(to);
        adjListTo.pushBack(&from);
    }
}

public const f<bool> Graph.hasCycles() {
    return false; // ToDo: Implement
}

public const f<bool> Graph.isDirected() {
    return this.directed;
}

public const f<bool> Graph.isDAG() {
    return this.directed && !this.hasCycles();
}

public const p Graph.toGraphviz(StringStream& ss) {
    const string graphType = this.directed ? "digraph" : "graph";
    const string edgeSep = this.directed ? "->" : "--";
    ss << graphType << " G {\n";

    // Emit all vertices
    foreach const Vertex<T>& v : this.vertices {
        ss << "  \"" << toString(v.value) << "\";\n";
    }

    // Emit all edges
    foreach const dyn pair : this.adjList {
        const T& srcValue = pair.getFirst().value;
        foreach const Vertex<T>* dst : pair.getSecond() {
            ss << "  \"" << toString(srcValue) << "\" " << edgeSep << " \"" << toString(dst.value) << "\";\n";
        }
    }

    ss << "}";
}
