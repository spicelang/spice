f<dyn> calledFunction(int mandatoryParam, dyn optionalParam = true) {
    printf("Mandatory: %d", mandatoryParam);
    printf("Optional: %d", optionalParam);

    /*string output = "";
    for int i = 0; i < 5; i++ {
        output += "test";
    }
    printf("Output: %s", output);*/

    return 0.1;
}

f<dyn> calledFunction(bool testBool) {
    printf("Bool: %d", testBool);
    return 0.3;
}

f<int> main() {
    dyn res = calledFunction(1, false);
    printf("Result: %d", res);
    calledFunction(false);
    return 0;
}