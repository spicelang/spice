import "std/data/vector";
import "std/io/filepath";
import "std/io/file";
import "std/text/transformation";

public type CSVRow interface {

}

type T int|double|string;
type RowType dyn;

public type CSVTable<RowType> struct {
    Vector<String> headers
    Vector<CSVRow> rows
}

/**
 * Parser for CSV files/strings.
 *
 * Usage:
 * ```spice
 * import "std/io/csv";
 * FilePath filePath = FilePath("path/to/file.csv");
 * CSVParser parser = CSVParser(filePath);
 * CSVTable table = parser.parse();
 * ```
 */
public type CSVParser<RowType> struct {
    CSVTable<RowType> table
    String input
    char separator
}

public p CSVParser.ctor(FilePath& csvFile, char separator = ',') {
    Result<String> fileContentOrError = readFile(csvFile.toString());
    this.input = fileContentOrError.unwrap();
    this.separator = separator;
}

public p CSVParser.ctor(const String& csvString, char separator = ',') {
    this.input = csvString;
    this.separator = separator;
}

public f<CSVTable<RowType>&> CSVParser.parse() {
    // Read the CSV file line by line
    Vector<String> lines = split(this.input, '\n');
    if (lines.isEmpty()) {
        return this.table;
    }
    // Parse the header line
    String headerLine = lines[0];
    Vector<String> headers = split(headerLine, this.separator);
    this.table.headers = headers;
    // Parse the data lines


    return this.table;
}
