import "std/io/dir" as dir;

f<int> main() {
    bool exists = dir.dirExists("./test");
    printf("Exists: %d\n", exists);
}