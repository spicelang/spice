p testProc(int t) {
    printf("%d", t);
}

f<int> main() {
    dyn test;
    testProc(test);
}