f<int> main() {
    int size = 5;
    int[size] array;
    printf("%d", sizeof(array));
}