import "std/data/vector";
import "std/text/print";
import "std/io/file" as io;

f<int> main() {
  dyn v = Vector<String>();
  v.pushBack(String("Hello"));
  v.pushBack(String("World!"));
  createFile("output.txt");
  const File file = openFile("output.txt", io::MODE_WRITE);

  for int i = 0; i < v.getSize(); i++ {
    String str = v.get(i);
    file.writeString((string) str.getRaw());
  }

  file.close();
}


/*type TestStruct struct {
    long lng
    String str
    int i
}

f<TestStruct> fct(int& ref) {
    TestStruct ts = TestStruct{ 6l, String("test string"), ref };
    return ts;
}

f<int> main() {
    int test = 987654;
    const TestStruct res = fct(test);
    printf("Long: %d\n", res.lng);
    printf("String: %s\n", res.str.getRaw());
    printf("Int: %d\n", res.i);
}*/