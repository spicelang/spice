/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec.Vector<pair.Pair<int, string>> pairVector = vec.Vector<pair.Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair.Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

f<int> main() {
    int[10][10] a;
    for int i = 0; i < 10; i++ {
        for int j = 0; j < 10; j++ {
            a[i][j] = i * j;
        }
    }
    printf("Cell [1,3]: %d", a[1][3]);
}