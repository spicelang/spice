const bool SIZE = false;

f<int> main() {
    short[SIZE] test;
}