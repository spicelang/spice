type Base struct {
    int x = 123
}

type A struct {
    compose Base base
    int a = 456
}

type B struct {
    compose Base base
    int b = 789
}

f<int> main() {
    unsafe {
        A a;
        Base* base = cast<Base*>(&a);
        B* b = cast<B*>(base);
        printf("b.b: %d\n", b.b);
    }
}