public type Any struct {
    bool test
}