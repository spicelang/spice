ext<byte*> malloc(long);

type ShoppingItem struct {
    string name
    double amount
    string unit
}

type ShoppingCart struct {
    string label
    ShoppingItem* items
}

f<ShoppingCart> newShoppingCart() {
    ShoppingItem* items;
    unsafe {
        items = (ShoppingItem*) malloc(sizeof(type ShoppingItem) * 3l);
        items[0] = ShoppingItem { "Spaghetti", 100.0, "g" };
        items[1] = ShoppingItem { "Rice", 125.5, "g" };
        items[2] = ShoppingItem { "Doughnut", 6.0, "pcs" };
    }
    return ShoppingCart { "Shopping Cart", items };
}

f<int> main() {
    ShoppingCart shoppingCart = newShoppingCart();
    unsafe {
        printf("Shopping cart item 1: %s\n", shoppingCart.items[1].name);
    }
}