// Imports
import "std/io/filepath";
import "std/io/file";
import "std/type/result";
import "../reader/code-loc";

public type Reader struct {
    File file
    string filename
    char curChar = '\0'
    bool moreToRead = true
    unsigned long line = 1l
    unsigned long col = 0l
}

public p Reader.ctor(const string inputFileName) {
    this.filename = inputFileName;
    Result<File> result = openFile(inputFileName, MODE_READ);
    this.file = result.unwrap();
    if !file.isOpen() {

    }
}

public p Reader.dtor() {
    file.close();
}

/**
 * @brief Get the previously read character
 *
 * @return char Last character
 */
public f<char> Reader.getChar() {
    return this.curChar;
}

/**
 * @brief Get the code location of the previously read character
 *
 * @return CodeLoc Code location
 */
public f<CodeLoc> Reader.getCodeLoc() {
    return CodeLoc(this.line, this.col, this.filename);
}

/**
 * @brief Advance the reader by one character
 */
public p Reader.advance() {
    assert !this.isEOF();
    if !this.file.get(this.curChar) {
        this.moreToRead = false;
    }
    if this.curChar == '\n' {
        this.line++;
        this.col = 0l;
    }
    this.col++;
}

/**
 * @brief Advance the reader by one character and check if this char equals the
 * expected
 *
 * @param c Expected char
 */
public p Reader.expect(char c) {
    assert this.curChar == c;
    this.advance();
}

/**
 * @brief Check if we are at the end of the input file
 *
 * @return At the end or not
 */
public f<bool> Reader.isEOF() {
    return !this.moreToRead;
}