f<int> main() {
    for dyn i = 0; i < 10; i+=2 {
        printf("Step %d\n", i);
    }
}

/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec::Vector<pair::Pair<int, string>> pairVector = vec.Vector<pair::Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair::Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

/*import "std/runtime/string_rt" as _rt_str;

f<int> main() {
    //_rt_str::String s = _rt_str::String("Test");
    //printf("%s", s.getRaw());
     // Plus
    printf("Result: %s\n", "Hello " + "World!");
    string s1 = "Hello " + "World!";
    printf("Result: %s\n", s1);
    // Mul
    printf("Result: %s\n", 4s * "Hi");
    string s2 = "Hello " * 5;
    printf("Result: %s\n", s2);
    printf("Result: %s\n", 20 * 'a');
    string s3 = 2 * 'c' * 7;
    printf("Result: %s\n", s3);
    //printf("%s", s1 + s2);
}*/

/*public f<int> src(int x, int y) {
    return x + (x | -x);
}

public f<int> tgt(int x) {
    return x & (x - 1);
}

f<int> main() {
    printf("Src: %d\n", src(21, 10));
    printf("Tgt: %d\n", tgt(21));
}*/