int GLOBAL_VARIABLE = 12;