import "std/type/result";
import "std/type/error";

// Constants
const unsigned long INITIAL_ALLOC_COUNT = 5l;
const unsigned int RESIZE_FACTOR = 2;

// Add generic type definition
type T dyn;

/**
 * A vector in Spice is a commonly used data structure, which can be used to represent a list of items.
 *
 * Time complexity:
 * Insert: O(1)
 * Delete: O(n * m); n = deleted elements, m = moved elements
 * Search: O(n)
 *
 * Vectors pre-allocate space using an initial size and a resize factor to not have to re-allocate
 * with every item pushed.
 */
public type Vector<T> struct {
    heap T* contents        // Pointer to the first data element
    unsigned long capacity  // Allocated number of items
    unsigned long size      // Current number of items
}

public p Vector.ctor(unsigned long initAllocItems = INITIAL_ALLOC_COUNT) {
    // Allocate space for the initial number of elements
    const long itemSize = sizeof(type T) / 8l;
    assert itemSize != 0l;
    unsafe {
        Result<heap byte*> allocResult = sAlloc(itemSize * initAllocItems);
        this.contents = (heap T*) allocResult.unwrap();
    }
    this.size = 0l;
    this.capacity = initAllocItems;
}

public p Vector.ctor(unsigned int initAllocItems) {
    this.ctor((long) initAllocItems);
}

public p Vector.ctor(unsigned long initAllocItems, const T& defaultValue) {
    // Allocate space for the initial number of elements
    this.ctor(initAllocItems);
    // Fill in the default values
    for int index = 0; index < initAllocItems; index++ {
        unsafe {
            this.contents[index] = defaultValue;
        }
    }
    this.size = initAllocItems;
}

/**
 * Checks if the vector contains any items at the moment
 *
 * @return Empty or not empty
 */
public f<bool> Vector.isEmpty() {
    return this.size == 0;
}

/**
 * Checks if the vector exhausts its capacity and needs to resize at the next call of push
 *
 * @return Full or not full
 */
public f<bool> Vector.isFull() {
    return this.size == this.capacity;
}

/**
 * Add an item at the end of the vector
 */
public p Vector.pushBack<T>(const T& item) {
    // Check if we need to re-allocate memory
    if this.isFull() {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Insert the element at the back
    unsafe {
        this.contents[(int) this.size++] = item;
    }
}

/**
 * Get an item at a certain index
 *
 * @return item at index
 */
public f<T&> Vector.get(unsigned long index) {
    if index >= this.size { panic(Error("Access index out of bounds")); }
    unsafe {
        return this.contents[index];
    }
}

/**
 * Get an item at a certain index
 *
 * @return item at index
 */
public f<T&> Vector.get(unsigned int index) {
    return this.get((unsigned long) index);
}

/**
 * Get the first item in the vector
 *
 * @return item at index 0
 */
public f<T&> Vector.front() {
    return this.get(0);
}

/**
 * Get the last item in the vector
 *
 * @return item at index size - 1
 */
public f<T&> Vector.back() {
    return this.get(this.size - 1);
}

/**
 * Removes all items from the vector
 */
public p Vector.clear() {
    this.size = 0l;
}

/**
 * Reserves `itemCount` items
 */
public p Vector.reserve(unsigned long itemCount) {
    if itemCount > this.capacity {
        this.resize(itemCount);
    }
}

/**
 * Reserves `itemCount` items
 */
public p Vector.reserve(unsigned int itemCount) {
    if itemCount > this.capacity {
        this.resize((long) itemCount);
    }
}

/**
 * Retrieve the current size of the vector
 *
 * @return Current size of the vector
 */
public f<long> Vector.getSize() {
    return this.size;
}

/**
 * Retrieve the current capacity of the vector
 *
 * @return Current capacity of the vector
 */
public f<long> Vector.getCapacity() {
    return this.capacity;
}

/**
 * Frees allocated memory that is not used by the queue
 */
public p Vector.pack() {
    // Return if no packing is required
    if this.isFull() { return; }
    // Pack the array
    this.resize(this.size);
}

public f<bool> operator==<T>(const Vector<T>& lhs, const Vector<T>& rhs) {
    // Compare the sizes
    if lhs.size != rhs.size { return false; }
    // Compare the contents
    for int index = 0; index < lhs.size; index++ {
        if lhs.contents[index] != rhs.contents[index] { return false; }
    }
    return true;
}

public f<bool> operator!=<T>(const Vector<T>& lhs, const Vector<T>& rhs) {
    return !(lhs == rhs);
}

/**
 * Re-allocates heap space for the queue contents
 */
p Vector.resize(unsigned long itemCount) {
    // Allocate the new memory
    const long itemSize = sizeof(type T) / 8l;
    assert itemSize != 0l;
    unsafe {
        heap byte* oldAddress = (heap byte*) this.contents;
        unsigned long newSize = (unsigned long) (itemSize * itemCount);
        Result<heap byte*> allocResult = sRealloc(oldAddress, newSize);
        this.contents = (heap T*) allocResult.unwrap();
    }
    // Set new capacity
    this.capacity = itemCount;
}