f<int> main() {
    int calcResult = "test" | 6;
    double otherResult = false & 6.7;
    string thirdResult = 6.7 ^ "test";
}