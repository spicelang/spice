f<int> main() {
    int new = 90;
    printf("New is: %s", new);
}