// Imports
import "bootstrap/reader/code-loc";

// Enums
public type TokenType enum {
    INVALID = 0,
    // Keyword tokens
    TYPE_DOUBLE = 1,
    TYPE_INT = 2,
    TYPE_SHORT = 3,
    TYPE_LONG = 4,
    TYPE_BYTE = 5,
    TYPE_CHAR = 6,
    TYPE_STRING = 7,
    TYPE_BOOL = 8,
    TYPE_DYN = 9,
    CONST = 10,
    SIGNED = 11,
    UNSIGNED = 12,
    INLINE = 13,
    PUBLIC = 14,
    HEAP = 15,
    COMPOSE = 16,
    F = 17,
    P = 18,
    IF = 19,
    ELSE = 20,
    SWITCH = 21,
    CASE = 22,
    DEFAULT = 23,
    ASSERT = 24,
    FOR = 25,
    FOREACH = 26,
    DO = 27,
    WHILE = 28,
    IMPORT = 29,
    BREAK = 30,
    CONTINUE = 31,
    FALLTHROUGH = 32,
    RETURN = 33,
    AS = 34,
    STRUCT = 35,
    INTERFACE = 36,
    TYPE = 37,
    ENUM = 38,
    OPERATOR = 39,
    ALIAS = 40,
    UNSAFE = 41,
    NIL = 42,
    MAIN = 43,
    PRINTF = 44,
    SIZEOF = 45,
    ALIGNOF = 46,
    LEN = 47,
    PANIC = 48,
    EXT = 49,
    CAST = 50,
    TRUE = 51,
    FALSE = 52,
    // Operator tokens
    LBRACE = 53,
    RBRACE = 54,
    LPAREN = 55,
    RPAREN = 56,
    LBRACKET = 57,
    RBRACKET = 58,
    LOGICAL_OR = 59,
    LOGICAL_AND = 60,
    BITWISE_OR = 61,
    BITWISE_XOR = 62,
    BITWISE_AND = 63,
    PLUS_PLUS = 64,
    MINUS_MINUS = 65,
    PLUS_EQUAL = 66,
    MINUS_EQUAL = 67,
    MUL_EQUAL = 68,
    DIV_EQUAL = 69,
    REM_EQUAL = 70,
    SHL_EQUAL = 71,
    SHR_EQUAL = 72,
    AND_EQUAL = 73,
    OR_EQUAL = 74,
    XOR_EQUAL = 75,
    PLUS = 76,
    MINUS = 77,
    MUL = 78,
    DIV = 79,
    REM = 80,
    NOT = 81,
    BITWISE_NOT = 82,
    GREATER = 83,
    LESS = 84,
    GREATER_EQUAL = 85,
    LESS_EQUAL = 86,
    SHL = 87,
    SHR = 88,
    EQUAL = 89,
    NOT_EQUAL = 90,
    ASSIGN = 91,
    QUESTION_MARK = 92,
    SEMICOLON = 93,
    COLON = 94,
    COMMA = 95,
    DOT = 96,
    ARROW = 97,
    SCOPE_ACCESS = 98,
    ELLIPSIS = 99,
    FCT_ATTR_PREAMBLE = 100,
    MOD_ATTR_PREAMBLE = 101,
    // Regex tokens
    DOUBLE_LIT = 102,
    INT_LIT = 103,
    SHORT_LIT = 104,
    LONG_LIT = 105,
    CHAR_LIT = 106,
    STRING_LIT = 107,
    IDENTIFIER = 108,
    TYPE_IDENTIFIER = 109,
    // Skipped tokens
    DOC_COMMENT = 110,
    BLOCK_COMMENT = 111,
    LINE_COMMENT = 112,
    EOF = 113
}

public type Token struct {
    public TokenType tokenType
    public String text
    public CodeLoc codeLoc
}

public p Token.ctor(TokenType tokenType) {
    this.tokenType = tokenType;
}

public p Token.ctor(TokenType tokenType, String text, const CodeLoc& codeLoc) {
    this.tokenType = tokenType;
    this.text = text;
    this.codeLoc = codeLoc;
}

public p Token.ctor(TokenType tokenType, string text, const CodeLoc& codeLoc) {
    this.ctor(tokenType, String(text), codeLoc);
}

public p Token.print() {
    printf("Token(type=%d, text=\"%s\", line=%d, col: %d)\n", this.tokenType, this.text, this.codeLoc.line, this.codeLoc.col);
}