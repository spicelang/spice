f<int> main() {
    int j;
    for j = 0; j < 5; j++ {
        printf("For round: %d", j);
    }
    return 0;
}