//import "std/runtime/string" as str;
//import "std/type/string" as tyStr;

f<int> main() {
    char a = 'a';
    byte a = 12;
    //string a = "Hello ";
    //string b = "World!";
    //printf("String a: %s\n", a);
    //printf("String b: %s\n", b);
    //printf("String a length: %d\n", tyStr.len(a));
    //printf("String a+b: %s", a + b);
}