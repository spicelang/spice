/*import "std/data/vector";
import "std/text/print";
import "std/io/file" as io;

f<int> main() {
  dyn v = Vector<String>();
  v.pushBack(String("Hello"));
  v.pushBack(String("World!"));
  createFile("output.txt");
  const File file = openFile("output.txt", io::MODE_WRITE);

  for int i = 0; i < v.getSize(); i++ {
    const String& str = v.get(i);
    file.writeString(str.getRaw());
  }

  file.close();
}*/

type intref struct {
    int test
}

f<bool> fn(const int& ref) {
    return false;
}

f<int> main() {
    const int x = 123;
    fn(x);
}