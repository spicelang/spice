// Std imports
import "std/data/map";
import "std/data/vector";

// Own imports
import "../ast/ast-nodes";
import "../symboltablebuilder/type";
import "../symboltablebuilder/symbol-table-entry";
import "../symboltablebuilder/type-specifiers";
import "../model/capture";
import "../model/generic-type";
import "../model/function";
import "../model/interface";

public type ScopeType enum {
    GLOBAL,
    FUNC_PROC_BODY,
    STRUCT,
    INTERFACE,
    ENUM,
    IF_ELSE_BODY,
    WHILE_BODY,
    FOR_BODY,
    FOREACH_BODY,
    SCOPE_THREAD_BODY,
    UNSAFE_BODY
}

/**
 * Class for storing information about symbols of the AST. Symbol tables are meant to be arranged in a tree structure,
 * so that you can navigate with the getParent() and getChild() methods up and down the tree.
 */
public type SymbolTable struct {
    SymbolTable* parent
    ScopeType scopeType
    Map<string, SymbolTable *> children
    Map<string, SymbolTableEntry> symbols
    Map<string, Capture> captures
    Map<string, GenericType> genericTypes
    Map<string, Map<string, Function>> functions // <code-loc, vector-of-representations>
    Map<string, Function*> functionAccessPointers
    Map<string, Map<string, Struct>> structs // <code-loc, vector-of-representations>
    Map<string, Struct*> structAccessPointers
    Map<string, Interface> interfaces

    bool inMainSourceFile
    bool isSourceFileRootScope
    bool isShadowTable
    bool capturingRequired
}

public p SymbolTable.ctor(
    const SymbolTable* parent,
    const ScopeType scopeType,
    const bool inMainSourceFile = false,
    const bool isSourceFileRoot = false
) {
    this.parent = parent;
    this.scopeType = scopeType;

    this.inMainSourceFile = inMainSourceFile;
    this.isSourceFileRootScope = isSourceFileRoot;
    this.isShadowTable = false;
    this.capturingRequired = false;
}

/**
 * Insert a new symbol into the current symbol table. If it is a parameter, append its name to the paramNames vector
 *
 * @param name Name of the symbol
 * @param symbolType Type of the symbol
 * @param specifiers Specifiers of the symbol
 * @param state State of the symbol (declared or initialized)
 * @param declNode AST node where the symbol is declared
 */
public p SymbolTable.insert(
    const string name,
    const Type symbolType,
    const TypeSpecifiers specifiers,
    const SymbolState state,
    const AstNode* declNode
) {
    bool global = this.parent == nil<SymbolTable*>;
    unsigned int orderIndex = this.symbols.getSize();
    // Insert into symbols map
    symbols.insert(SymbolTableEntry{name, symbolType, this, specifiers, state, declNode, orderIndex, global});
}

/**
 * Insert a new anonymous symbol into the current symbol table.
 * The anonymous symbol will be identified via the definition code location
 *
 * @param symbolType Type of the symbol
 * @param declNode AST node where the symbol is declared
 */
public p SymbolTable.insertAnonymous(const Type symbolType, const AstNode* declNode) {
    string name = "anon." + declNode.codeLoc.toString();
    this.insert(name, symbolType, TypeSpecifiers(symbolType), SymbolState.DECLARED, declNode);
    this.lookupAnonymous(declNode.codeLoc).used = true;
}

/**
 * Check if a symbol exists in the current or any parent scope and return it if possible
 *
 * @param name Name of the desired symbol
 * @return Desired symbol / nullptr if the symbol was not found
 */
public f<SymbolTableEntry*> SymbolTable.lookup(const string name) {
    // Check if the symbol exists in the current scope. If yes, take it
    SymbolTableEntry* entry = this.lookupStrict(name);
    if entry != nil<SymbolTableEntry*> { // Symbol was not found in the current scope
        // We reached the root scope, the symbol does not exist at all
        if parent == nil<SymbolTable*> { return nil<SymbolTableEntry*>; }
        // If there is a parent scope, continue the search there
        entry = this.parent.lookup(name);
        // Symbol was also not found in all the parent scopes, return nullptr
        if entry == nil<SymbolTable*> { return nil<SymbolTableEntry*>; }

        // Check if this scope requires capturing and capture the variable if appropriate
        if this.capturingRequired && !this.captures.contains(name) && !entry.ty.isOneOf({TY_IMPORT, TYPE_FUNCTION, TY_PROCEDURE}) {
            this.captures.insert(name, Capture(entry));
        }
    }
    return entry;
}

/**
 * Check if a symbol exists in the current scope and return it if possible
 *
 * @param name Name of the desired symbol
 * @return Desired symbol / nullptr if the symbol was not found
 */
public f<SymbolTableEntry*> SymbolTable.lookupStrict(const string name) {
    if name.isEmpty() { return nil<SymbolTableEntry*>; }
    // Check if a symbol with this name exists in this scope
    if this.symbols.contains(name) { return &this.symbols.get(name); }
    // Check if a capture with this name exists in this scope
    if this.captures.contains(name) { return &this.captures.get(name).capturedEntry; }
    // Otherwise, return a nullptr
    return nil<SymbolTableEntry*>;
}

/**
 * Check if an order index exists in the current or any parent scope and returns it if possible.
 * Warning: Unlike the `lookup` method, this one doesn't consider the parent scopes
 *
 * @param orderIndex Order index of the desired symbol
 * @return Desired symbol / nullptr if the symbol was not found
 */
public f<SymbolTableEntry*> SymbolTable.lookupStrictByIndex(const unsigned int orderIndex) {
    // ToDo
    return nil<SymbolTableEntry*>;
}

/**
 * Check if a global variable exists in any of the imported modules and return it if found
 *
 * @param globalName Name of the global variable
 * @param skipThisScope Skip the current scope while searching
 * @return Desired symbol / nullptr if the global was not found
 */
public f<SymbolTableEntry*> SymbolTable.lookupGlobal(const string globalName, const bool skipThisScope = false) {
    // Search in the current scope
    if !skipThisScope {
        SymbolTableEntry* globalSymbol = this.lookupStrict(globalName);
        if globalSymbol != nil<SymbolTableEntry*> { return globalSymbol; }
    }
    // Loop through all children to find the global var
    // ToDo
    return nil<SymbolTableEntry*>;
}

/**
 * Check if an anonymous symbol exists in the current scope and return it if possible
 *
 * @param codeLoc Definition code loc
 * @return Anonymous symbol
 */
public f<SymbolTableEntry*> SymbolTable.lookupAnonymous(const CodeLoc codeLoc) {
    return this.lookup("anon." + codeLoc.toString());
}

/**
 * Check if a capture exists in the current or any parent scope scope and return it if possible
 *
 * @param captureName Name of the desired captured symbol
 * @return Capture / nullptr if the capture was not found
 */
public f<Capture> SymbolTable.lookupCapture(const string captureName) {
    // Check if the capture exists in the current scope. If yes, take it
    Capture* capture = this.lookupCaptureStrict(name);
    if capture != nil<Capture*> { return capture; }

    // We reached the root scope, the symbol does not exist at all
    if this.parent == nil<SymbolTable*> { return nullptr; }

    return this.parent.lookupCapture(name);
}

/**
 * Check if a capture exists in the current scope and return it if possible
 *
 * @param captureName Name of the desired captured symbol
 * @return Capture / nullptr if the capture was not found
 */
public f<Capture> SymbolTable.lookupCaptureStrict(const string captureName) {

}

/**
 * Search for a symbol table by its name, where a function is defined. Used for function calls to function/procedures
 * which were linked in from other modules
 *
 * @param tableName Name of the desired table
 * @return Desired symbol table
 */
public f<SymbolTable*> SymbolTable.lookupTable(const string tableName) {
    // If not available in the current scope, search in the parent scope
    if !this.children.contains(tableName) {
        return this.parent != nil<SymbolTable*> ? this.parent.lookupTable(tableName) : nil<SymbolTable*>;
    }
    // Otherwise, return the entry
    return this.children.get(tableName);
}

/**
 * Create a child leaf for the tree of symbol tables and return it
 *
 * @param childBlockName Name of the child scope
 * @param type Type of the child scope
 * @return Newly created child table
 */
public f<SymbolTable*> SymbolTable.createChildBlock(const string tableName, const ScopeType scopeType) {
    // ToDo
}

/**
 * Insert a new generic type in this scope
 *
 * @param typeName Name of the generic type
 * @param genericType Generic type itself
 */
public p SymbolTable.insertGenericType(const string typeName, const GenericType genericType) {
    this.genericTypes.insert(typeName, genericType);
}

/**
 * Search for a generic type by its name. If it was not found, the parent scopes will be searched.
 * If the generic type does not exist at all, the function will return a nullptr.
 *
 * @param typeName Name of the generic type
 * @return Generic type
 */
public f<GenericType> SymbolTable.lookupGenericType(const string typeName) {
    if this.genericTypes.contains(typeName) {
        return &this.genericTypes.get(typeName);
    }
    return this.parent != nil<SymbolTable*> ? this.parent.lookupGenericType(typeName) : nil<GenericType*>;
}

/**
 * Mount in symbol tables manually. This is used to hook in symbol tables of imported modules into the symbol table of
 * the source file, which imported the modules
 *
 * @param childBlockName Name of the child block
 * @param childBlock Child symbol table
 * @param alterParent Set the current symbol table as parent of the mounted one
 */
public p SymbolTable.mountChildBlock(const string childBlockName, const SymbolTable *childBlock, const bool alterParent = true) {
    if alterParent {
        childBlock.parent = this;
    }
    this.children.insert(childBlockName, childBlock);
}

/**
 * Rename the scope of a symbol table. This is useful for realizing function overloading by storing a function with not
 * only its name, but also its signature
 *
 * @param oldName Old name of the child table
 * @param newName New name of the child table
 */
public p SymbolTable.renameChildBlock(const string oldName, const string newName) {
    // ToDo
}

/**
 * Duplicates the child block by copying it. The duplicated symbols point to the original ones.
 *
 * @param oldName Original name of the child block
 * @param newName New block name
 */
public p SymbolTable.copyChildBlock(const string oldName, const string newName) {
    assert this.children.contains(oldName);
    SymbolTable* originalChildBlock = this.children.get(oldName);
    // Copy child block
    // ToDo
    // Save the new child block
    this.children.insert(newName, newChildBlock);
}

/**
 * Navigate to a child table of the current one in the tree structure
 *
 * @param tableName Name of the child table
 * @return Pointer to the child symbol table
 */
public f<SymbolTable*> SymbolTable.getChild(const string tableName) {
    if this.children.isEmpty() || !this.children.contains(tableName) { return nil<SymbolTable*>; }
    return children.get(tableName);
}

/**
 * Retrieve all variables that can be freed, because the ref count went down to 0.
 *
 * @param filterForDtorStructs Get only struct variables
 * @return Variables that can be de-allocated
 */
public f<Vector<SymbolTableEntry*>> SymbolTable.getVarsGoingOutOfScope(const bool filterForDtorStructs = false) {
    assert this.parent != nil<SymbolTable*>; // Should not be called in root scope
    Vector<SymbolTableEntry*> varsGoingOutOfScope;

    // Collect all variables in this scope
    // ToDo

    // Collect all variables in the child scopes
    // ToDo

    return varsGoingOutOfScope;
}

/**
 * Returns all symbols of the current table
 *
 * @return Map of names and the corresponding symbol table entries
 */
public f<Map<string, SymbolTableEntry>*> SymbolTable.getSymbols() {
    return &this.symbols;
}

/**
 * Returns all captures of the current table
 *
 * @return Map of names and the corresponding capture
 */
public f<Map<string, Capture>*> SymbolTable.getCaptures() {
    return &this.captures;
}

/**
 * Get the number of fields if this is a struct scope
 *
 * @return Number of fields
 */
public f<long> SymbolTable.getFieldCount() {
    assert this.scopeType == ScopeType.STRUCT;
    unsigned long fieldCount = 0l;
    // ToDo
    return fieldCount;
}

/**
 * Insert a function object into this symbol table scope
 *
 * @param function Function object
 * @param err Error factory
 */
public f<Function*> SymbolTable.insertFunction(const Function *function) {
    const AstNode *declNode = function.declNode;
    // ToDo
    return nil<Function*>;
}

/**
 * Check if there is a function in this scope, fulfilling all given requirements and if found, return it.
 * If more than one function matches the requirement, an error gets thrown
 *
 * @param currentScope Current scope
 * @param callFunctionName Function name requirement
 * @param callThisType This type requirement
 * @param callArgTypes Argument types requirement
 * @param node Declaration node for a potential error message
 * @return Matched function or nullptr
 */
public f<Function*> SymbolTable.matchFunction(
    SymbolTable* currentScope,
    const string callFunctionName,
    const Type callThisType,
    const Vector<Type>* callArgTypes,
    const AstNode* node
) {
    Vector<Function*> matches;

    // Loop through functions and add any matches to the matches vector
    // ToDo

    if matches.isEmpty() { return nil<Function*>; }

    // Throw error if more than one function matches the criteria
    if matches.getSize() > 1 {
        // ToDo
    }

    // Add function access pointer for function call
    if currentScope != nil<SymbolTable*> {
        string suffix = callFunctionName == DTOR_FUNCTION_NAME ? callFunctionName : "";
        currentScope.insertFunctionAccessPointer(matches.front(), node.codeLoc, suffix);
    }

    return matches.front();
}

/**
 * Retrieve the manifestations of the function, defined at defToken
 *
 * @param defCodeLoc Definition code location
 * @return Function manifestations
 */
public f<Map<string, Function>*> SymbolTable.getFunctionManifestations(const CodeLoc defCodeLoc) {
    string codeLocStr = defCodeLoc.toString();
    return this.functions.contains(codeLocStr) ? this.functions.get(codeLocStr) : nil<Map<string, Function>*>;
}

/**
 * Add function access pointer to the current scope
 *
 * @param spiceFunc Function
 * @param codeLoc Call code location
 * @param suffix Key suffix
 */
public p SymbolTable.insertFunctionAccessPointer(
    const Function* spiceFunc,
    const CodeLoc codeLoc,
    const string suffix
) {
    string mapKey = codeLoc.toString() + ":" + suffix;
    this.functionAccessPointers.insert(mapKey, spiceFunc);
}

/**
 * Get the function access pointer by code location
 *
 * @param codeLoc Code location
 * @param suffix Key suffix
 *
 * @return Function pointer for the function access
 */
public f<Function*> SymbolTable.getFunctionAccessPointer(const CodeLoc codeLoc, const string suffix) {
    string mapKey = codeLoc.toString() + ":" + suffix;
    return this.functionAccessPointers.contains(mapKey) ? this.functionAccessPointers.get(mapKey) : nil<Function*>;
}

/**
 * Insert a substantiated function into the function list. If the list already contains a function with the same signature,
 * an exception will be thrown
 *
 * @param function Substantiated function
 * @param declNode Declaration AST node
 */
f<Function*> SymbolTable.insertSubstantiatedFunction(const Function spiceFunc, const AstNode* declNode) {
    // ToDo
}

/**
 * Insert a struct object into this symbol table scope
 *
 * @param spiceStruct Struct object
 */
public f<Struct*> SymbolTable.insertStruct(const Struct *spiceStruct) {
    // Open a new struct declaration pointer list. Which gets filled by the 'insertSubstantiatedStruct' method
    string codeLocStr = spiceStruct.declNode.codeLoc.toString();
    //this.stucts.insert(codeLocStr, );
    return this.insertSubstantiatedStruct(spiceStruct, spiceStruct.declNode);
}

/**
 * Check if there is a struct in this scope, fulfilling all given requirements and if found, return it.
 * If more than one struct matches the requirement, an error gets thrown
 *
 * @param currentScope Current scope
 * @param structName Struct name
 * @param templateTypes Template type requirements
 * @param node Declaration node for the error message
 * @return Matched struct or nullptr
 */
public f<Struct*> SymbolTable.matchStruct(
    SymbolTable* currentScope,
    const string structName,
    const Vector<Type>* templateTypes,
    const AstNode* node
) {
    Vector<Struct*> matches;

    // ToDo
}

/**
 * Retrieve the manifestations of the struct, defined at defToken
 *
 * @return Struct manifestations
 */
public f<Map<string, Struct>*> SymbolTable.getStructManifestations(const CodeLoc defCodeLoc) {
    string codeLocStr = defCodeLoc.toString();
    if !this.structs.contains(codeLocStr) {
        // ToDo
    }
    return this.structs.get(codeLocStr);
}

/**
 * Add struct access pointer to the current scope
 *
 * @param codeLoc Reference code location
 * @param struct Struct
 */
public p SymbolTable.insertStructAccessPointer(const CodeLoc codeLoc, const Struct* spiceStruct) {
    this.structAccessPointers.insert(codeLoc.toString, spiceStruct);
}

/**
 * Get the next struct access in order of visiting
 *
 * @return Struct pointer for the struct access
 */
public f<Struct*> SymbolTable.getStructAccessPointer(const CodeLoc codeLoc, const string suffix = "") {
    string codeLocStr = codeLoc.toString();
    if !this.structAccessPointers.contains(codeLocStr) {
        // ToDo
    }
    return this.structAccessPointers.get(codeLocStr);
}

/**
 * Insert a substantiated struct into the struct list. If the list already contains a struct with the same signature,
 * an exception will be thrown
 *
 * @param s Substantiated struct
 * @param declNode Declaration AST node
 */
f<Struct*> SymbolTable.insertSubstantiatedStruct(const Struct spiceStruct, const AstNode* declNode) {
    // ToDo
}

/**
 * Retrieve an interface instance by its name
 *
 * @param interfaceName Name of the interface
 * @return Interface object
 */
public f<Interface*> SymbolTable.lookupInterface(const string interfaceName) {
    if !this.interfaces.contains(interfaceName) { return nil<Interface*>; }
    return &this.interfaces.get(interfaceName);
}

/**
 * Insert an interface object into this symbol table scope
 *
 * @param i Interface object
 */
public p SymbolTable.insertInterface(const Interface* i) {
    // Add interface to interface list
    assert !this.interfaces.contains(i.name);
    this.interfaces.insert(i.name, i);
    // Add symbol table entry for the interface
    this.insert(i.name, Type(TY_INTERFACE), i.specifiers, INITIALIZED, i.declNode);
}

/**
 * Retrieves compiler warnings from this table
 */
public f<Vector<CompilerWarning>> SymbolTable.collectWarnings() {
    // ToDo
}

/**
 * Checks if this symbol table is imported
 *
 * @param askingScope Symbol table, which asks whether the current one is imported from its point of view or not
 *
 * @return Imported / not imported
 */
public f<bool> SymbolTable.isImportedBy(const SymbolTable* askingScope) {
    // ToDo
}