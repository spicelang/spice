f<int> main() {
    string food = "Pizza";
    string* ptr = &food;

    printf("Pointer address: %p, value: %s", ptr, *ptr);

    *ptr = "Burger";

    dyn restoredFood = *ptr;
    printf("Restored value: %s", restoredFood);

    printf("Restored value address: %p\n", &restoredFood);
}