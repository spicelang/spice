f<int> main() {
    // Simple address check
    int test = 123;
    int& testRef = test;
    assert &test == &testRef;

    // Try operators
    testRef += 12;
    assert test == 135;
    testRef -= 11;
    assert test == 124;
    testRef = 123;
    assert test == 123;
    testRef = testRef + 4;
    assert test == 127;
    testRef = testRef - 4;
    assert test == 123;

    printf("All assertions passed!");
}

/*import "std/iterator/number-iterator";

f<int> main() {
    foreach long idx, short item : range(1s, 19s) {
        printf("%d: %d\n", idx, item);
    }

    printf("All assertions passed!");
}*/