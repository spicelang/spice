/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/net/socket" as socket;

f<int> main() {
    socket.Socket s = socket.openServerSocket(8080s, 2);
    printf("Error code: %d", s.errorCode);
    //s.close();
}*/



import "std/time/delay" as delay;
import "std/os/system" as sys;

f<int> main() {
    printf("Starting threads ...\n");
    //int coreCount = sys.getCPUCoreCount() / 2;
    for int i = 1; i <= 7; i++ {
        printf("Starting thread %d ...\n", i);
        thread {
            printf("Tid: %d, i: %d\n", tid(), i);
        }
    }
    delay.delay(3000);
    printf("Hello from original\n");
}