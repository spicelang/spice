f<int> main() {
    /*printf("Array1:\n");
    short arraySize1 = 3s;
    int[arraySize1] array1 = {1, 2, 3};
    foreach dyn item : array1 {
        printf("Item: %d\n", item);
    }

    printf("\nArray2:\n");
    long arraySize2 = 2l;
    string[arraySize2] array2;
    array2[0] = "one";
    array2[1] = "two";
    foreach dyn item : array2 {
        printf("Item: %s\n", item);
    }

    printf("\nArray3:\n");
    int arraySize3 = 3;
    int[arraySize3] array3 = {1, arraySize3, arraySize3};
    foreach dyn item : array3 {
        printf("Item: %d\n", item);
    }*/

    printf("\nArray4:\n");
    int arraySize4 = 3;
    int[arraySize4] array4;
    array4 = {1, arraySize4, arraySize4};
    foreach dyn item : array4 {
        printf("Item: %d\n", item);
    }
}