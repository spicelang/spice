import "std/io/cli-parser";

type CliOptions struct {
    bool sayHi = false
}

p callback(bool& value) {
    printf("Callback called with value %d\n", value);
}

f<int> main(int argc, string[] argv) {
    CliParser parser = CliParser("Test Program", "This is a simple test program");
    parser.setVersion("v0.1.0");
    parser.setFooter("Copyright (c) Marc Auberer 2021-2023");

    CliOptions options;
    parser.addFlag("--hi", options.sayHi, "Say hi to the user");
    parser.addFlag("--callback", callback, "Call a callback function");
    parser.addFlag("-cb", p(bool& value) {
        printf("CB called with value %d\n", value);
    }, "Call a callback function");

    parser.parse(argc, argv);

    // Print hi if requested
    if options.sayHi {
        printf("Hi!\n");
    }
}

/*import "std/os/thread-pool";

f<int> main() {
    ThreadPool tp = ThreadPool(3s);
    tp.enqueue(p() {
        printf("Hello from task 1\n");
    });
    tp.enqueue(p() {
        printf("Hello from task 2\n");
    });
    tp.enqueue(p() {
        printf("Hello from task 3\n");
    });
    tp.enqueue(p() {
        printf("Hello from task 4\n");
    });
}*/

/*type T int|long;

type TestStruct<T> struct {
    T _f1
    unsigned long length
}

p TestStruct.ctor(const unsigned long initialLength) {
    this.length = initialLength;
}

p TestStruct.printLength() {
    printf("%d\n", this.length);
}

type Alias alias TestStruct<long>;

f<int> main() {
    Alias a = Alias{12345l, (unsigned long) 54321l};
    a.printLength();
    dyn b = Alias(12l);
    b.printLength();
}*/

/*type TestStruct struct {
    long lng
    String str
    int i
}

p TestStruct.dtor() {}

f<TestStruct> fct(int& ref) {
    TestStruct ts = TestStruct{ 6l, String("test string"), ref };
    return ts;
}

f<int> main() {
    int test = 987654;
    const TestStruct res = fct(test);
    printf("Long: %d\n", res.lng);
    printf("String: %s\n", res.str.getRaw());
    printf("Int: %d\n", res.i);
}*/