type T int|double;

public type Vector<T> struct {
    public T data
}

public p Vector.setData<T>(T data) {
    this.data = data;
    foreach int item : reverse(items) {

    }
}