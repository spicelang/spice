/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

f<int> main() {
    int[7] intArray = { 1, 5, 4, 0, 12, 12345, 9 };
    /*foreach (int index, int item : intArray) {
        printf("Item for index %d, %d", index, item);
    }*/
    foreach (const int idx = 2, const int item : intArray) {
        printf("Item for index %d, %d", idx, item);
        idx++;
    }
    /*foreach const int item : intArray {
        printf("Item: %d", idx);
        printf("Item: %d", item);
    }*/
}