f<int> main() {
    int[5] array = { 1, 2, 3, 4, 5 };
    foreach double item : array {
        printf("Item: %f", item);
    }
}