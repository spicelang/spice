type Test struct {
    int i = 5.67
}

f<int> main() {}