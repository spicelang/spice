#![core.compiler.alwaysKeepOnNameCollision = true]

// Link external functions
ext f<heap byte*> malloc(unsigned long);
ext f<heap byte*> realloc(heap byte*, unsigned long);
ext p free(heap byte*);
ext p memcpy(heap byte*, heap byte*, unsigned long);
ext f<int> memcmp(const heap byte*, const heap byte*, unsigned long);

// Generic type defs
type T dyn;

/**
  * Allocates a new block of memory of the given size.
  *
  * @param size The size of the block to allocate.
  * @return A pointer to the allocated block, or an error if the allocation failed.
  */
public f<Result<heap byte*>> sAlloc(unsigned long size) {
    heap byte* ptr = malloc(size);
    return ptr != nil<heap byte*> ? ok(ptr) : err<heap byte*>("OOM occurred in sAlloc!");
}

/**
  * Allocates a new block of memory of the given size.
  * This panics in case of an out of memory situation.
  *
  * @param size The size of the block to allocate.
  * @return A pointer to the allocated block
  */
public f<heap byte*> sAllocUnsafe(unsigned long size) {
    heap byte* ptr = malloc(size);
    if ptr != nil<heap byte*> { return ptr; }
    panic(Error("OOM occurred in sAllocUnsafe!"));
}

/**
  * Reallocates a block of memory to the given size.
  * Subsequently moves the data from the old memory space to the new one.
  *
  * @param ptr The pointer to the block to reallocate.
  * @param size The new size of the block.
  * @return A pointer to the reallocated block, or an error if the reallocation failed.
  */
public f<Result<heap byte*>> sRealloc(heap byte* ptr, unsigned long size) {
    if ptr == nil<heap byte*> { return err<heap byte*>("Original pointer is nil!"); }
    if size == 0l { return err<heap byte*>("Size is 0!"); }
    heap byte* newPtr = realloc(ptr, size);
    return newPtr != nil<heap byte*> ? ok(newPtr) : err<heap byte*>("OOM occurred in sRealloc!");
}

/**
  * Reallocates a block of memory to the given size.
  * Subsequently moves the data from the old memory space to the new one.
  * This panics in case of invalid input or an out of memory situation.
  *
  * @param ptr The pointer to the block to reallocate.
  * @param size The new size of the block.
  * @return A pointer to the reallocated block, or an error if the reallocation failed.
  */
public f<heap byte*> sReallocUnsafe(heap byte* ptr, unsigned long size) {
    if ptr == nil<heap byte*> { panic(Error("Original pointer is nil!")); }
    if size == 0l { panic(Error("Size is 0!")); }
    heap byte* newPtr = realloc(ptr, size);
    if newPtr == nil<heap byte*> {
        panic(Error("OOM occurred in sReallocUnsafe!"));
    }
    return newPtr;
}

/**
  * Copies a block of memory to a new block of memory.
  *
  * @param oldPtr The pointer to the block to copy.
  * @param newPtr The pointer to the new block to copy to.
  * @param size The size of the block to copy.
  * @return A pointer to the copied block, or an error if the copy failed.
  */
public f<Result<heap byte*>> sCopy(heap byte* oldPtr, heap byte* newPtr, unsigned long size) {
    if oldPtr == nil<heap byte*> | newPtr == nil<heap byte*> {
        return err<heap byte*>("Cannot copy from or to nil pointer!");
    }
    memcpy(newPtr, oldPtr, size);
    return ok(newPtr);
}

/**
  * Copies a block of memory to a new block of memory.
  *
  * @param oldPtr The pointer to the block to copy.
  * @param newPtr The pointer to the new block to copy to.
  * @param size The size of the block to copy.
  * @return A pointer to the copied block, or an error if the copy failed.
  */
public f<heap byte*> sCopyUnsafe(heap byte* oldPtr, heap byte* newPtr, unsigned long size) {
    if oldPtr == nil<heap byte*> | newPtr == nil<heap byte*> {
        panic(Error("Cannot copy from or to nil pointer!"));
    }
    memcpy(newPtr, oldPtr, size);
    return newPtr;
}

/**
  * Moves the ownership of a heap pointer from oldPtr to the return value.
  * After this operation, oldPtr is set to nil to prevent double frees.
  *
  * @param oldPtr The pointer to move ownership from
  * @return The moved pointer
  */
public f<heap T*> sMove<T>(heap T*& oldPtr) {
    result = oldPtr;
    oldPtr = nil<heap T*>;
}

/**
 * Allocates memory for a new instance of the given type on the heap.
 * Note: This function panics if the allocation fails.
 *
 * @return A pointer to the heap-allocated instance
 */
public f<heap T*> sNew<T>() {
    unsafe {
        // Allocate memory for the instance
        Result<heap byte*> res = sAlloc(sizeof<T>());
        return cast<heap T*>(res.unwrap());
    }
}

/**
 * Allocates memory for a new instance of the given type on the heap.
 * Note: This function panics if the allocation fails.
 *
 * @param val The value to put into the heap-allocated memory
 * @return A pointer to the heap-allocated instance
 */
public f<heap T*> sNew<T>(const T& val) {
    unsafe {
        // Allocate memory for the instance
        Result<heap byte*> res = sAlloc(sizeof<T>());
        result = cast<heap T*>(res.unwrap());
        // Copy the value into the heap-allocated memory
        sCopy(cast<heap byte*>(&val), cast<heap byte*>(result), sizeof<T>());
    }
}

/**
 * Allocates memory for a new instance of the given type on the heap.
 *
 * @param ptr The pointer to the heap-allocated memory
 * @param val The value to put into the heap-allocated memory
 * @return A pointer to the heap-allocated instance
 */
public f<T*> sPlacementNew<T>(heap byte* ptr, const T& val) {
    unsafe {
        // Copy the value into the heap-allocated memory
        sCopy(cast<heap byte*>(&val), ptr, sizeof<T>());
        return cast<T*>(ptr);
    }
}

/**
 * Destroys the given object by calling its dtor if available
 *
 * @param obj The object to destroy
 */
public p sDestruct<T>(T& obj) {
    obj.dtor();
}

/**
  * Frees a block of memory.
  * The pointer is zeroed out after freeing the memory to prevent accidental double frees.
  *
  * @param ptr The pointer to the block to free.
  */
public p sDealloc(heap byte*& ptr) {
    if ptr == nil<heap byte*> { return; }
    free(ptr);
    ptr = nil<heap byte*>; // Zero out to prevent accidental double frees
}

/**
 * Destroys the given heap-allocated instance and frees the memory.
 *
 * @param ptr The pointer to the heap-allocated instance
 */
public p sDelete<T>(heap T*& ptr) {
    sDestruct(*ptr);
    unsafe {
        sDealloc(cast<heap byte*&>(ptr));
    }
}

/**
 * Yields the ownership of the given heap pointer.
 * After this operation, the original pointer is set to nil to prevent double frees.
 *
 * @param ptr The pointer to yield ownership from
 * @return The yielded pointer
 */
public f<T*> sYieldOwnership<T>(heap T*& ptr) {
    result = ptr;
    ptr = nil<heap T*>;
}

/**
 * Compares the memory behind pointer A and pointer B for equality.
 *
 * @param a Pointer A
 * @param b Pointer B
 * @return Is memory equal
 */
public f<bool> sCompare<T>(const heap T* a, const heap T* b, unsigned long size) {
    unsafe {
        return memcmp(cast<const byte*>(a), cast<const byte*>(b), size) == 0;
    }
}
