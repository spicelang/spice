public type IGenericType interface {

}
