f<int> main() {
    int[10] testArray = { 1, 2, 3, 4, 5, 6, 7, 8, 9, 10};
    printf("Test: %d\n", testArray[15]);
}