// External declarations
ext f<long> strtol(string, char**, int);

// Converts a string to a double
public f<double> toDouble(string input) {
    // ToDo: implement
    return 0.0;
}

// Converts a string to an int
public f<int> toInt(string input, int base = 10) {
    return (int) toLong(input, base);
}

// Converts a string to a short
public f<short> toShort(string input, int base = 10) {
    return (short) toLong(input, base);
}

// Converts a string to a long
public f<long> toLong(string input, int base = 10) {
    char* endPtr = nil<char*>;
    result = strtol(input, &endPtr, base);
    // Check if the conversion was successful
    if (((string) endPtr) == input || *endPtr != '\0') { return 0l; }
}

// Converts a string to a byte
public f<byte> toByte(string input, int base = 10) {
    return (byte) ((int) toLong(input, base));
}

// Converts a string to a char
public f<char> toChar(string input) {
    return input[0];
}

// Converts a string to a bool
public f<bool> toBool(string input) {
    return input == "true";
}