ext<int> usleep(int);

f<int> main() {
    printf("Starting one thread ...\n");
    thread {
        usleep(500 * 1000);
        printf("Hello from the thread 1\n");
    }
    thread {
        usleep(200 * 1000);
        printf("Hello from the thread 2\n");
    }
    usleep(1000 * 1000);
    printf("Hello from original\n");
}

/*const int THREAD_COUNT = 8;

f<int> fib(int n) {
    if n <= 2 { return 1; }
    return fib(n - 1) + fib(n - 2);
}

f<int> main() {
    byte*[THREAD_COUNT] threads = {};
    for unsigned int i = 0; i < THREAD_COUNT; i++ {
        threads[i] = thread {
            printf("Thread returned with result: %d\n", fib(46));
        };
        printf("%p\n", threads[i]);
    }
    printf("Started all threads. Waiting for results ...\n");
    join(threads);
    printf("Program finished");
}*/