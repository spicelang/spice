#![core.compiler.alwaysKeepOnNameCollision = true]

import "std/iterator/array-iterator";

// Generic type definitions
type I dyn; // Item type

/**
 * Convenience wrapper for creating a simple array iterator
 */
public inline f<ArrayIterator<I>> iterate<I>(I[] array, unsigned long size) {
    return ArrayIterator<I>(array, size);
}