import "std/data/optional";

f<int> main() {
    Optional<int> iO = Optional<int>(12);
    printf("%d", iO.get());
}