type T dyn;
type TRes dyn;

// -------------------------------------- cast<T>(x) --------------------------------------

p castInner<TRes, T>(T lhs, TRes expectedResult) {
    const TRes actualResult = cast<TRes>(lhs);
    assert actualResult == expectedResult;
}

p castInnerUnsafe<TRes, T>(T lhs, TRes expectedResult) {
    unsafe {
        const TRes actualResult = cast<TRes>(lhs);
        assert actualResult == expectedResult;
    }
}

p castTest() {
    // Identity casts
    castInner<double, double>(1.123, 1.123);
    castInner<int, int>(123, 123);
    castInner<short, short>(3457s, 3457s);
    castInner<long, long>(23068763214l, 23068763214l);
    castInner<byte, byte>(cast<byte>(324), cast<byte>(324));
    castInner<char, char>('+', '+');
    castInner<string, string>("test", "test");
    castInner<bool, bool>(true, true);
    bool b = false;
    castInner<bool*, bool*>(&b, &b);
    // Lhs double
    castInner<double, int>(1, 1.0);
    castInner<double, short>(1s, 1.0);
    castInner<double, long>(1l, 1.0);
    // Lhs int
    castInner<int, double>(1.0, 1);
    castInner<int, short>(1s, 1);
    castInner<int, long>(1l, 1);
    castInner<int, byte>(cast<byte>(1), 1);
    castInner<int, char>('A', 65);
    // Lhs short
    castInner<short, double>(1.0, 1s);
    castInner<short, int>(1, 1s);
    castInner<short, long>(1l, 1s);
    // Lhs long
    castInner<long, double>(1.0, 1l);
    castInner<long, int>(1, 1l);
    castInner<long, short>(1s, 1l);
    // Lhs byte
    castInner<byte, int>(56, cast<byte>(56));
    castInner<byte, char>('8', cast<byte>(56));
    // Lhs char
    castInner<char, int>(57, '9');
    castInner<char, short>(57s, '9');
    castInner<char, long>(57l, '9');
    castInner<char, byte>(cast<byte>(57), '9');
    // Special casts
    // cast<const char*>(string)
    String str = String("test");
    castInner<string, const char*>(cast<const char*>(str.getRaw()), "test");
    // cast<char[]>(string)
    castInner<string, const char[]>(['t', 'e', 's', 't', '\0'], "test");
    // cast<string>(const char*)
    castInner<const char*, string>("test", cast<const char*>(str.getRaw()));
    // cast<any*>(any*)
    castInnerUnsafe<int*, short*>(nil<short*>, nil<int*>);
}

f<int> main() {
    castTest(); // cast<T>(x)
    printf("All assertions passed!");
}