f<int> main() {
    short s = (short) 10;
    s++;
    long l = (long) 10;
    printf("Short: %d, Long: %d\n", s, l);
}