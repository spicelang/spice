/**
 * Returns a formatted storage string (e.g. 1.4 MB for 1,500,000)
 *
 * @return Formatted size string
 */
public f<string> formatStorageSize(long bytes) {
    // ToDo when string concatenation works
    return "";
}

/**
 * Returns the given text in caps
 *
 * @return Text in caps
 */
public f<string> toUpper(string text) {
    const char shiftOffset = (char) 32;
    const char min = (char) 97;
    const char max = (char) 122;

    foreach char c : text {
        if c >= min && c <= max {
            c += shiftOffset;
        }
    }
    return text;
}

/**
 * Returns the given text in all-lower letters
 *
 * @return Text in all-lower letters
 */
public f<string> toLower(string text) {
    const char shiftOffset = (char) 32;
    const char min = (char) 65;
    const char max = (char) 90;

    foreach char c : text {
        if c >= min && c <= max {
            c -= shiftOffset;
        }
    }
    return text;
}

/**
 * Returns the given text in capitalized form
 *
 * @return Capitalized text
 */
public f<string> capitalize(string text) {
    if text[0] >= (char) 97 && text[0] <= (char) 122 {
        text[0] += (char) 32;
    }
    return text;
}