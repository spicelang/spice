import "std/test/lifetime-object";

f<LifetimeObject> spawnLO() {
    return LifetimeObject();
}

f<int> main() {
    // Ignored return value of ctor
    printf("Ignored return value of ctor:\n");
    {
        LifetimeObject();
    }

    // Normal lifecycle
    printf("Normal lifecycle:\n");
    {
        LifetimeObject lo = LifetimeObject(); // ctor call
        LifetimeObject loCopy = lo; // copy ctor call
    } // dtor calls for both lo and loCopy at end of scope

    // Return from lambda as value
    printf("Return from lambda as value:\n");
    {
        const f<LifetimeObject>() spawnLO = f<LifetimeObject>() {
            return LifetimeObject();
        };

        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    // Return from lambda as reference
    printf("Return from lambda as reference:\n");
    {
        LifetimeObject loOrig = LifetimeObject();
        const f<LifetimeObject&>() spawnLO = f<LifetimeObject&>() {
            return loOrig;
        };

        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    // Return from lambda as const reference
    printf("Return from lambda as const reference:\n");
    {
        LifetimeObject loOrig = LifetimeObject();
        const f<const LifetimeObject&>() spawnLO = f<const LifetimeObject&>() {
            return loOrig;
        };

        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    // Return from function as value
    printf("Return from function as value:\n");
    {
        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }
}