// Std imports
import "std/text/stringstream";

// Own imports
import "bootstrap/reader/code-loc";

public type CompilerWarningType enum {
    UNUSED_FUNCTION,
    UNUSED_PROCEDURE,
    UNUSED_METHOD,
    UNUSED_STRUCT,
    UNUSED_INTERFACE,
    UNUSED_IMPORT,
    UNUSED_FIELD,
    UNUSED_ENUM_ITEM,
    UNUSED_ALIAS,
    UNUSED_VARIABLE,
    UNUSED_RETURN_VALUE,
    UNREACHABLE_CODE,
    SHADOWED_VARIABLE,
    IDENTITY_CAST,
    SINGLE_GENERIC_TYPE_CONDITION,
    BOOL_ASSIGN_AS_CONDITION,
    ASYNC_LAMBDA_CAPTURE_RULE_VIOLATION,
    UNINSTALL_FAILED,
    VERIFIER_DISABLED
}

/**
 * Compiler warning template engine
 */
public type CompilerWarning struct {
    String warningMessage
}

/**
 * Constructor: Used in case that the exact code position where the warning occurred is known
 *
 * @param codeLoc Code location, where the warning occurred
 * @param warningType Type of the warning
 * @param message Warning message suffix
 */
public p CompilerWarning.ctor(const CodeLoc& codeLoc, const CompilerWarningType warningType, const string message) {
    StringStream msg;
    msg << "[Warning] " << codeLoc.toPrettyString() << ": " << this.getMessagePrefix(warningType) << ": " << message;
    this.warningMessage = msg.str();
}

/**
 * Constructor: Used in case the exact code position where the warning occurred is not known
 *
 * @param warningType Type of the warning
 * @param message Warning message suffix
 */
public p CompilerWarning.ctor(const CompilerWarningType warningType, const string message) {
    StringStream msg;
    msg << "[Warning] " << this.getMessagePrefix(warningType) << ": " << message;
    this.warningMessage = msg.str();
}

/**
 * Print the compiler warning to the standard error output
 */
public p CompilerWarning.print() {
    printf("%s", this.warningMessage);
}

/**
 * Get the prefix of the warning message for a particular error
 *
 * @param type Type of the warning
 * @return Prefix string for the warning type
 */
f<string> CompilerWarning.getMessagePrefix(const CompilerWarningType warningType) {
    switch warningType {
        case CompilerWarningType::UNUSED_FUNCTION: { return "Unused function"; }
        case CompilerWarningType::UNUSED_PROCEDURE: { return "Unused procedure"; }
        case CompilerWarningType::UNUSED_METHOD: { return "Unused method"; }
        case CompilerWarningType::UNUSED_STRUCT: { return "Unused struct"; }
        case CompilerWarningType::UNUSED_INTERFACE: { return "Unused interface"; }
        case CompilerWarningType::UNUSED_IMPORT: { return "Unused import"; }
        case CompilerWarningType::UNUSED_FIELD: { return "Unused field"; }
        case CompilerWarningType::UNUSED_ENUM_ITEM: { return "Unused enum item"; }
        case CompilerWarningType::UNUSED_ALIAS: { return "Unused type alias"; }
        case CompilerWarningType::UNUSED_VARIABLE: { return "Unused variable"; }
        case CompilerWarningType::UNUSED_RETURN_VALUE: { return "Unused return value"; }
        case CompilerWarningType::UNREACHABLE_CODE: { return "Unreachable code detected"; }
        case CompilerWarningType::SHADOWED_VARIABLE: { return "Shadowed variable"; }
        case CompilerWarningType::IDENTITY_CAST: { return "Identity cast"; }
        case CompilerWarningType::SINGLE_GENERIC_TYPE_CONDITION: { return "Only one type condition"; }
        case CompilerWarningType::BOOL_ASSIGN_AS_CONDITION: { return "Bool assignment as condition"; }
        case CompilerWarningType::ASYNC_LAMBDA_CAPTURE_RULE_VIOLATION: { return "Lambda violates async lambda capture rule"; }
        case CompilerWarningType::UNINSTALL_FAILED: { return "Uninstall failed"; }
        case CompilerWarningType::VERIFIER_DISABLED: { return "Verifier disabled"; }
        default: { panic(Error("Unknown warning")); }
    }
}