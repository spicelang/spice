import "std/io/file";

f<int> main() {
    string filename = "./test-file.txt";
    bool _ = deleteFile(filename); // Ensure that the file is not present in the beginning

    assert !fileExists(filename);
    assert createFile(filename);
    assert fileExists(filename);
    assert deleteFile(filename);
    assert !fileExists(filename);

    printf("All assertions passed!");
}