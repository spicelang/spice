import "os-test2" as os;

f<int> main() {
    Vec test = Vec{1, false};
    test.print();
    return 0;
}