f<int> main() {
    long l = 1234l;
    long* lPtr = &l;
    int* iPtr;
    unsafe {
        iPtr = (int*) lPtr;
    }
    printf("Int: %d\n", *iPtr);
}