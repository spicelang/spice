f<int> main() {
    (1) = 4;
}