import "std/type/bool" as boolTy;

f<int> main() {
    printf("Result: %d\n", boolTy.toInt(true));
}