type Visitor struct {

}

type SymbolTable struct {

}

type Visitable interface {
    f<bool> accept(Visitor*)
}

type AstNode struct : Visitable {

}

type AstEntryNode struct : Visitable {
    AstNode astNode
    SymbolTable* fctScope
    bool hasArgs
}

f<int> main() {
    dyn entryNode = AstEntryNode{};
    printf("%d", entryNode.hasArgs);
}

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

/*public f<bool> src(bool x, bool y) {
    return ((x ? 1 : 4) & (y ? 1 : 4)) == 0;
}

public f<int> tgt(int x, int y) {
    return x ^ y;
}

f<int> main() {
    printf("Result: %d, %d", src(false, true), tgt(0, 1));
}*/