type TestStruct struct {
    long a
    short b
    string a
}

f<int> main() {}