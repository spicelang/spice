// Imports
import "std/text/print";
import "std/os/cmd";
import "std/io/cli-parser";

/**
 * Representation of the various cli options
 */
public type CliOptions struct {
    public String mainSourceFile // e.g. main.spice
    public String targetTriple   // In format: <arch><sub>-<vendor>-<sys>-<abi>
    public String targetArch
    public String targetVendor
    public String targetOs
    public bool execute
    public bool isNativeTarget
    public String cacheDir
    public String outputDir      // Where the object files go. Should always be a temp directory
    public String outputPath     // Where the output binary goes.
    public unsigned short compileJobCount // O for auto
    public bool ignoreCache
    public bool printDebugOutput
    public bool dumpCST
    public bool dumpAST
    public bool dumpIR
    public bool dumpAssembly
    public bool dumpSymbolTables
    public bool disableAstOpt
    public short optLevel // -O0 = 0, -O1 = 1, -O2 = 2, -O3 = 3, -Os = 4, -Oz = 5
    public bool generateDebugInfo
    public bool disableVerifier
    public bool testMode
}

/**
 * Helper class to setup the cli interface and command line parser
 */
public type CliInterface struct {
    CliParser cliParser
    public CliOptions cliOptions
    public bool shouldCompile
    public bool shouldInstall
    public bool shouldExecute
}

public p CliInterface.ctor() {
    // Initialize cli object
    this.cliOptions = CliOptions{
        /* mainSourceFile */ String(""),
        /* targetTriple */ String(""),
        /* targetArch */ String(""),
        /* targetVendor */ String(""),
        /* targetOs */ String(""),
        /* execute */ false,
        /* isNativeTarget */ false,
        /* cacheDir */ String(""),
        /* outputDir */ String(""),
        /* outputPath */ String(""),
        /* compileJobCount */ 0s,
        /* ignoreCache */ false,
        /* printDebugOutput */ false,
        /* dumpCST */ false,
        /* dumpAST */ false,
        /* dumpIR */ false,
        /* dumpAssembly */ false,
        /* dumpSymbolTables */ false,
        /* disableAstOpt */ false,
        /* optLevel */ 2s,
        /* generateDebugInfo */ false,
        /* disableVerifier */ false,
        /* testMode */ false
    };
    this.shouldCompile = false;
    this.shouldInstall = false;
    this.shouldExecute = false;
}

public p CliInterface.createInterface() {
    this.cliParser = CliParser("Spice", "Spice programming language");
    this.cliParser.setFooter("Copyright (c) Marc Auberer 2021-2023");

    // Add version flag
    this.cliParser.setVersion("Spice version 0.14.3\nbuilt by: GitHub Actions\n\n(c) Marc Auberer 2021-2023");

    // Create sub-commands
    this.addBuildSubcommand();
    this.addRunSubcommand();
    this.addInstallSubcommand();
    this.addUninstallSubcommand();

    // ToDo: extend
}

/**
 * Validates if all necessary cli options were provided.
 *
 * @throws InvalidCliOptionsException if there were an invalid combination of cli options provided
 */
public p CliInterface.validate() {
    if ((this.cliOptions.targetArch.isEmpty() && this.cliOptions.targetVendor.isEmpty() && this.cliOptions.targetOs.isEmpty()) ||
        (!this.cliOptions.targetArch.isEmpty() && !this.cliOptions.targetVendor.isEmpty() && !this.cliOptions.targetOs.isEmpty())) {
        // ToDo: throw cli error
    }

    // Error out when opt level > 0 and debug info enabled
    if (this.cliOptions.optLevel > 0 && this.cliOptions.generateDebugInfo) {
        // ToDo: throw cli error
    }
}

/**
 * Initialize the cli options based on the input of the user
 */
public p CliInterface.enrich() {
    // Propagate target information
    if this.cliOptions.targetTriple.isEmpty() && this.cliOptions.targetArch.isEmpty() {
        // ToDo: Extend
    }

    // Dump AST, IR and symbol table if all debug output is enabled
    if this.cliOptions.printDebugOutput {
        this.cliOptions.dumpAST = true;
        this.cliOptions.dumpIR = true;
        this.cliOptions.dumpSymbolTables = true;
    }
}

/**
 * Add build subcommand to cli interface
 */
p CliInterface.addBuildSubcommand() {
    // Create sub-command itself
    // ToDo: Extend
}

/**
 * Add run subcommand to cli interface
 */
p CliInterface.addRunSubcommand() {
    // Create sub-command itself
    // ToDo: Extend
}

/**
 * Add install subcommand to cli interface
 */
p CliInterface.addInstallSubcommand() {
    // Create sub-command itself
    // ToDo: Extend
}

/**
 * Add uninstall subcommand to cli interface
 */
p CliInterface.addUninstallSubcommand() {
    // Create sub-command itself
    // ToDo: Extend
}

/**
 * Start the parsing process
 *
 * @param argc Argument count
 * @param argv Argument vector
 * @return Return code
 */
public f<int> CliInterface.parse(int argc, string[] argv) {
    return this.cliParser.parse(argc, argv);
}

/**
 * Executes the built executable
 */
p CliInterface.runBinary() {
    // Print status message
    if this.cliOptions.printDebugOutput {
        println("Running executable ...\n");
    }

    // Run executable
    execCmd(this.cliOptions.outputPath.getRaw());
}