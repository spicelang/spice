const int testInt = 0;
double testDouble = 1.5;
string testString = "";
bool testBool = true;
dyn testAuto = false;

// This is a test comment
f<int> testFunction(double doubleParam) {
    dyn number;
    number = 123;
    result = number | 5;

    while testDouble < 2.5 {
        for int i = 12; i < 15; i+=2 {
            result = 12;
        }
        testDouble += 2.0;
    }
}

p testProcedure(string stringParam, bool boolParam = false) {
    /* Test
    block
    comment */
    double result = testString == "" || testBool ? 5.0 : 1.4;
    if result == 5.0 { result = 3.0; }
    int result1 = testFunction(3.0);
    testProcedure("test", false);
}

f<int> main() {
    testProcedure();
    return 0;
}