type Visitor struct {}

type SymbolTable struct {}

type Visitable interface {
    f<bool> accept(Visitor*)
}

type AstNode struct : Visitable {}

type AstEntryNode struct : Visitable {
    AstNode astNode
    SymbolTable* fctScope
    bool hasArgs
}

f<int> main() {
    dyn entryNode = AstEntryNode{};
    printf("%d", entryNode.hasArgs);
}