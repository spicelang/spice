import "std/data/vector";
import "std/data/linked-list";
import "std/data/pair";
import "std/math/hash";

// Generic types for key and value
type K dyn;
type V dyn;

public type HashTable<K, V> struct {
    Vector<LinkedList<Pair<K, V>>> table
    unsigned long bucketCount
}

public p HashTable.ctor(unsigned long bucketCount = 100l) {
    this.bucketCount = bucketCount;
    this.table = Vector<LinkedList<Pair<K, V>>>(bucketCount);
}

public p HashTable.insert(const K& key, const V& value) {
    const unsigned long index = this.hash(key);
    LinkedList<Pair<K, V>>& bucket = this.table.get(index);
    foreach Pair<K, V>& pair : bucket.getIterator() {
        if pair.getFirst() == key {
            pair.setSecond(value);
            return;
        }
    }
    this.table.pushBack(LinkedList<Pair<K, V>>());
    LinkedList<Pair<K, V>>& bucket = this.table.back();
    bucket.pushBack(Pair<K, V>(key, value));
}

public p HashTable.delete(const K& key) {
    const unsigned long index = this.hash(key);
    const LinkedList<Pair<K, V>>& bucket = this.table.at(index);

    for unsigned long i = 0l; i < bucket.getSize(); i++ {
        Pair<K, V>& candidate = bucket.at(i);
        if candidate.getFirst() == key {
            bucket.remove(i);
            return;
        }
    }
}

public f<V*> HashTable.get(const K& key) {
    unsigned long index = this.hash(key);
    const LinkedList<Pair<K, V>>& bucket = this.table.at(index);

    for unsigned long i = 0l; i < bucket.getSize(); i++ {
        Pair<K, V>& candidate = bucket.at(i);
        if candidate.getFirst() == key {
            return &candidate.getSecond();
        }
    }
    return nil<V*>;
}

inline f<unsigned long> HashTable.hash(const K& key) {
    return hash(key) % this.bucketCount;
}