type TestStruct struct {
    unsigned int field1
    long field2
}

f<int> main() {
    int[9] intArray = {};
    printf("%d\n", sizeof(intArray));

    printf("%d\n", sizeof("Hello World!"));
}