// Generic types
type T dyn;

/**
 * Optionals in Spice are wrappers around values, that allow them to be empty.
 * This can be used as better alternative to nil for empty values.
 */
public type Optional<T> struct {
    T data
    bool isPresent = false
}

/**
 * Initialize optional without a value
 */
public p Optional.ctor() {}

/**
 * Initialize optional with an initial value
 *
 * @param data Initial data value
 */
public p Optional.ctor(const T& data) {
    this.data = data;
    this.isPresent = true;
}

/**
 * Set the value of the optional
 *
 * @param data New data value
 */
public inline p Optional.set(const T& data) {
    this.data = data;
    this.isPresent = true;
}

/**
 * Get the value of the optional
 *
 * @return Data value
 */
public inline f<T&> Optional.get() {
    if !this.isPresent { panic(Error("Optional payload is not present")); }
    return this.data;
}

/**
 * Get the value of the optional. If the optional is not present, return the default value
 *
 * @return Data value or default value
 */
public inline f<T&> Optional.orElse(T& defaultValue) {
    return this.isPresent ? this.data : defaultValue;
}

/**
  * Get the value of the optional. If the optional is not present, return the value of `getFct`
  *
  * @return Data value or value of the function
  */
public inline f<T&> Optional.orElseGet(f<T&>() getFct) {
    return this.isPresent ? this.data : getFct();
}

/**
 * Clears the value of the optional
 */
public inline p Optional.clear() {
    this.isPresent = false;
}

/**
 * Checks if a value is present at the moment
 *
 * @return Present or not
 */
public inline f<bool> Optional.isPresent() {
    return this.isPresent;
}

public f<bool> operator==<T>(const Optional<T>& lhs, const Optional<T>& rhs) {
    return lhs.isPresent == rhs.isPresent && lhs.data == rhs.data;
}

public f<bool> operator!=<T>(const Optional<T>& lhs, const Optional<T>& rhs) {
    return !(lhs == rhs);
}