// Imports
import "../lexer/token";