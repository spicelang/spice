import "source2";

f<int> add(int a, int b) {
    return a + b;
}

#[test]
f<bool> testAdd1() {
    assert add(1, 2) == 3;
    assert add(2, 2) == 4;
    assert add(3, 2) == 5;
    return true;
}

#[test]
f<bool> testAdd2() {
    assert add(5, -4) == 1;
    assert add(2, 8) == 10;
    assert add(-3, 5) == 2;
    return false;
}