/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/data/vector" as vector;

f<int> main() {
    dyn v = vector.Vector<int>{};
    v.push(4);
    v.push(2);
}*/

import "std/data/vector" as vec;

f<int> main() {
    dyn v1 = vec.Vector<int>{};
    //v1.ctor();
    //v1.pushBack(123);
    //v1.pushBack(90);
    //v1.dtor();
}