public f<int> functionInModuleB(int x, int y) {
  return x + y;
}