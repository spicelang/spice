import "std/text/print" as print;

type Test struct {
    int field1
    double field2
}

f<Test> Test.get() {
    printf("%d\n", this.field1);
    return *this;
}

p Test.print(bool b) {
    if b {
        printf("Content: %d, %f", this.field1, this.field2);
    }
}

f<int> main() {
    Test test = new Test { 5, 4.567 };
    dyn field1 = test.get().field1;
    printf("Field1: %d\n", field1);
    print.println("Test");
    printf("%d\n", test.field1);
    test.print(true);
}