type Test struct {
    int test
}

f<int> main() {
    Test t = Test{ 12 };
    printf("Test: %d", t.test);
}