#[test]
f<string> test() {
  return "failed";
}

f<int> main() {}