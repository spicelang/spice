f<int> main() {
    printf("Hello World!");
    return 0;
}