// Generic types
type T dyn;

public type Optional<T> struct {
    T data
    bool isPresent
}

public p Optional.ctor() {
    this.isPresent = false;
}

public p Optional.ctor(const T& data) {
    this.data = data;
    this.isPresent = true;
}

public inline p Optional.set(const T& data) {
    this.data = data;
    this.isPresent = true;
}

public inline f<T&> Optional.get() {
    return this.data;
}

public inline p Optional.clear() {
    this.isPresent = false;
}

public inline f<bool> Optional.isPresent() {
    return this.isPresent;
}