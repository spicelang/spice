import "std/data/vector" as v;

f<int> main() {
    dyn doubleVec = v.Vector<double>(3, 6.4);
    printf("Test: %f\n", doubleVec.get(0));
    printf("Test: %f\n", doubleVec.get(1));
    printf("Test: %f\n", doubleVec.get(2));
    printf("Test: %f\n", doubleVec.get(3));
    doubleVec.dtor();
}