const int COUNT;

f<int> main() {
    printf("Test");
}