import "std/math/fct" as fct;

f<int> main() {
    printf("Abs (int): %d\n", fct.abs(123));
    printf("Abs (int): %d\n", fct.abs(-137));
    printf("Abs (short): %d\n", fct.abs(56s));
    printf("Abs (short): %d\n", fct.abs(-3s));
    printf("Abs (long): %d\n", fct.abs(1234567890l));
    printf("Abs (long): %d\n", fct.abs(-987654321l));
    printf("Abs (double): %f\n", fct.abs(56.123));
    printf("Abs (double): %f\n", fct.abs(-348.12));

    printf("Floor (int): %d\n", fct.floor<int>(-348.12));
    long fl = fct.floor<long>(-348.12);
    printf("Floor (long): %d\n", fl);
    printf("Floor (short): %d\n", fct.floor<short>(-348.12));

    printf("Sin (double): %f\n", fct.sin(78.345));
    printf("Sin (int): %f\n", fct.sin(23));
    printf("Sin (short): %f\n", fct.sin(-68s));
    printf("Sin (long): %f\n", fct.sin(359l));

    printf("Cos (double): %f\n", fct.cos(78.345));
    printf("Cos (int): %f\n", fct.cos(23));
    printf("Cos (short): %f\n", fct.cos(-68s));
    printf("Cos (long): %f\n", fct.cos(359l));
}

/*type Visitor struct {

}

type SymbolTable struct {

}

type VisitableNode interface {
    f<bool> accept(Visitor*)
}

type AstNode struct : VisitableNode {

}

f<bool> AstNode.accept(Visitor* v) {
    return true;
}

type AstEntryNode struct : VisitableNode {
    AstNode astNode
    SymbolTable* fctScope
    bool hasArgs
}

f<bool> AstEntryNode.accept(Visitor* v) {
    return true;
}

f<int> main() {
    dyn entryNode = AstEntryNode{};
    printf("%d", entryNode.hasArgs);
}*/

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

/*public f<bool> src(bool x, bool y) {
    return ((x ? 1 : 4) & (y ? 1 : 4)) == 0;
}

public f<int> tgt(int x, int y) {
    return x ^ y;
}

f<int> main() {
    printf("Result: %d, %d", src(false, true), tgt(0, 1));
}*/