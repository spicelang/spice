f<int> main() {
    if 7 {
        printf("Test");
    }
}