public const int SIZE = 64;
public const long MIN_VALUE = -9223372036854775808;
public const long MAX_VALUE = 9223372036854775807;

// Converts a long to a double
public f<double> toDouble(long input) {
    return 0.0 + input;
}

// Converts a long to an int
public f<int> toInt(long input) {
    return (int) input;
}

// Converts a long to a short
public f<short> toShort(long input) {
    return (short) input;
}

// Converts a long to a byte
public f<byte> toByte(long input) {
    return (byte) input;
}

// Converts a long to a char
public f<char> toChar(long input) {
    return (char) input;
}

// Converts a long to a string
public f<string> toString(long input) {
    // ToDo: Implement (See https://github.com/golang/go/blob/master/src/strconv/itoa.go)
    return "";
}

// Converts a long to a boolean
public f<bool> toBool(long input) {
    return input >= 1;
}