f<int> main() {
    while true {
        break 0;
    }
}