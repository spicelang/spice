import "std/type/result";

// Link external functions
ext f<heap byte*> malloc(long);
ext f<heap byte*> realloc(heap byte*, int);
ext p free(heap byte*);
ext p memcpy(heap byte*, heap byte*, long);

/**
  * Allocates a new block of memory of the given size.
  *
  * @param size The size of the block to allocate.
  * @return A pointer to the allocated block, or an error if the allocation failed.
  */
public f<Result<heap byte*>> alloc(long size) {
    heap byte* ptr = malloc(size);
    return ptr != nil<heap byte*> ? ptr : err(nil<heap byte*>, "Out of memory occurred!");
}

/**
  * Reallocates a block of memory to the given size.
  *
  * @param ptr The pointer to the block to reallocate.
  * @param size The new size of the block.
  * @return A pointer to the reallocated block, or an error if the reallocation failed.
  */
public f<Result<heap byte*>> realloc(heap byte* ptr, long size) {
    heap byte* newPtr = realloc(ptr, size);
    return newPtr != nil<heap byte*> ? newPtr : err(nil<heap byte*>, "Out of memory occurred!");
}

/**
  * Copies a block of memory to a new block of memory.
  *
  * @param ptr The pointer to the block to copy.
  * @param size The size of the block to copy.
  * @return A pointer to the copied block, or an error if the copy failed.
  */
public f<Result<heap byte*>> copy(heap byte* ptr, long size) {
    heap byte* newPtr = malloc(size);
    if newPtr == nil<heap byte*> {
        return err(nil<heap byte*>, "Out of memory occurred!");
    }
    memcpy(newPtr, ptr, size);
    return newPtr;
}

/**
  * Frees a block of memory.
  * The pointer is zeroed out after freeing the memory to prevent accidental double frees.
  *
  * @param ptr The pointer to the block to free.
  */
public p dealloc(heap byte*& ptr) {
    free(ptr);
    ptr = nil<heap byte*>; // Zero out to prevent accidental double frees
}