import "std/type/bool" as Bool;

f<int> main() {
    printf("Result: %d", Bool.toInt(true));
}