f<int> main() {
    printf("%d", 6.23456);
}