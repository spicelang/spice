f<int> main() {
    long l = 1234l;
    long* lPtr = &l;
    int* iPtr = cast<int*>(lPtr);
    printf("Int: %d\n", *iPtr);
}