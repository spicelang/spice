import "std/type/char";

f<int> main() {
    // toDouble()
    double asDouble = toDouble('d');
    assert asDouble == 100.0;

    // toInt()
    int asInt = toInt('T');
    assert asInt == 84;

    // toShort()
    short asShort = toShort('j');
    assert asShort == 106s;

    // toLong()
    long asLong = toLong('K');
    assert asLong == 75l;

    // toString()
    String asString = toString('v');
    assert asString.getRaw() == "v";

    // toBool()
    bool asBool1 = toBool('1');
    assert asBool1 == true;
    bool asBool2 = toBool('0');
    assert asBool2 == false;

    printf("All assertions succeeded");
}