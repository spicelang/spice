#![core.linker.flag = "-pthread"]

// Type definitions
type Pthread_t alias long;
type Pthread_attr_t struct {
    unsigned byte detached
    char *ss_sp
    unsigned long ss_size
}

// Link external functions
ext f<int> pthread_create(Pthread_t* /*thread*/, Pthread_attr_t* /*attr*/, p() /*start_routine*/, byte* /*arg*/);
ext f<int> pthread_join(Pthread_t /*thread*/, byte** /*retval*/);
ext f<Pthread_t> pthread_self();

/**
 * Lightweight thread, that uses posix threads (pthread) under the hood.
 */
public type Thread struct {
    Pthread_t threadId
}

public p Thread.ctor(p() threadRoutine) {
    pthread_create(&this.threadId, nil<Pthread_attr_t*>, threadRoutine, nil<byte*>);
}

/**
 * Wait synchronous until the thread has terminated
 */
public p Thread.join() {
    pthread_join(this.threadId, nil<byte**>);
}

/**
 * Retrieve the ID of the current thread
 */
public f<Pthread_t> Thread.getId() {
    return this.threadId;
}

/**
 * Retrieve the ID of the current thread
 */
public f<Pthread_t> getThreadId() {
    return pthread_self();
}