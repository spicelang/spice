ext<int> usleep(int);

f<int> main() {
    printf("Starting threads ...\n");
    int capturedVariable = 0;
    for int i = 1; i <= 8; i++ { // Start 8 threads
        printf("Starting thread %d ...\n", i);
        thread {
            usleep(100 * i * 1000);
            capturedVariable *= 2;
            printf("Hello from the thread\n");
        }
    }
    usleep(1000 * 1000);
    printf("Hello from original\n");
}