import "test/functions" as functions;

f<int> main() {
    if true {
        printf("If");
    } else if false {
        printf("Else if");
    } else {
        printf("Else");
    }
    printf("Test\n");
}