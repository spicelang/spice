// Std imports
import "std/text/print";
import "std/os/cmd";
import "std/os/os";
import "std/os/filesystem";
import "std/io/cli-parser";
import "std/io/cli-subcommand";
import "std/io/cli-option";
import "std/io/filepath";
import "std/io/file";
import "std/time/time";
import "std/type/long";

// Own imports
import "util/common-util";
import "util/file-util";
import "util/compiler-warning";

// Constants
public const string TARGET_UNKNOWN = "unknown";
public const string TARGET_WASM32 = "wasm32";
public const string TARGET_WASM64 = "wasm64";
public const string ENV_VAR_DOCKERIZED = "SPICE_DOCKERIZED";

public type OptLevel enum {
    O0 = 0, // No optimization
    O1 = 1, // Only basic optimizations
    O2 = 2, // Default optimization level
    O3 = 3, // Aggressively optimize for performance
    Os = 4, // Optimize for code size
    Oz = 5  // Aggressively optimize for code size
}

public type BuildMode enum {
    DEBUG = 0,   // Default build mode, uses -O0 per default
    RELEASE = 1, // Build without debug information and with -O2 per default
    TEST = 2     // Build with test main function and always emit assertions
}
const string BUILD_MODE_DEBUG = "debug";
const string BUILD_MODE_RELEASE = "release";
const string BUILD_MODE_TEST = "test";

public type DumpSettings struct {
    public bool dumpCST = false
    public bool dumpAST = false
    public bool dumpSymbolTable = false
    public bool dumpTypes = false
    public bool dumpIR = false
    public bool dumpAssembly = false
    public bool dumpObjectFile = false
    public bool dumpToFiles = false
    public bool abortAfterDump = false
}

/**
 * Representation of the various cli options
 */
public type CliOptions struct {
    public FilePath mainSourceFile // e.g. main.spice
    public String targetTriple   // In format: <arch><sub>-<vendor>-<sys>-<abi>
    public String targetArch = String(TARGET_UNKNOWN)
    public String targetVendor = String(TARGET_UNKNOWN)
    public String targetOs = String(TARGET_UNKNOWN)
    public bool isNativeTarget = true
    public bool useCPUFeatures = true
    public bool execute = false
    public FilePath cacheDir                      // Where the cache files go. Should always be a temp directory
    public FilePath outputDir = FilePath("./")    // Where the object files go. Should always be a temp directory
    public FilePath outputPath                    // Where the output binary goes.
    public BuildMode buildMode = BuildMode::DEBUG // Default build mode is debug
    public unsigned int compileJobCount = 0       // O for auto
    public bool ignoreCache = false
    public String llvmArgs
    public bool printDebugOutput = false
    public DumpSettings dumpSettings
    public bool namesForIRValues = false
    public bool useLifetimeMarkers = false
    public OptLevel optLevel = OptLevel::O0 // Default optimization level for debug build mode is O0
    public bool useLTO = false
    public bool noEntryFct = false
    public bool generateTestMain = false
    public bool staticLinking = false
    public bool generateDebugInfo = false
    public bool disableVerifier = false
    public bool testMode = false
}

/**
 * Helper class to setup the cli interface and command line parser
 */
public type Driver struct {
    public CliOptions cliOptions
    public bool shouldCompile = false
    public bool shouldInstall = false
    public bool shouldUninstall = false
    public bool shouldExecute = false
    public bool dryRun = false // For unit testing purposes
    CliParser cliParser
}

public p Driver.init() {
    this.cliParser = CliParser("Spice", "Spice programming language");
    this.cliParser.setFooter("(c) Marc Auberer 2021-2025");

    // Add version flag
    this.cliParser.setVersion(buildVersionInfo());

    // Create sub-commands
    this.addBuildSubcommand();
    this.addRunSubcommand();
    this.addTestSubcommand();
    this.addInstallSubcommand();
    this.addUninstallSubcommand();

    // ToDo: Here we have a problem with passing the cautres. Curently the capture struct is stack-allocated. This stack
    // allocation goes out of scope at the end of the function, but used afterwards.
    /*this.cliParser.setRootCallback(p() {
        if this.shouldInstall || this.shouldUninstall {
            // Prepare the installation path
            FilePath installPath = getSpiceBinDir();
            installPath /= this.cliOptions.mainSourceFile.getBaseName();
            if !this.dryRun {
                // ToDo
            }

            // If the binary should be installed, set the output path to the Spice bin directory
            if this.shouldInstall {
                this.cliOptions.outputPath = installPath;
            }

            // If the binary should be uninstalled, check if the executable exists and uninstall it
            if this.shouldUninstall && !this.dryRun {
                if installPath.exists() && deleteFile(installPath.toString()) {
                    println("Successfully uninstalled");
                } else {
                    CompilerWarning warning = CompilerWarning(CompilerWarningType::UNINSTALL_FAILED, "The executable was not found at the expected location");
                    warning.print();
                }
            }
        }

        // Abort here if we do not need to compile
        if !this.shouldCompile {
            return;
        }

        // Set output path and dir
        if this.shouldExecute {
            this.cliOptions.execute = true;
            const long millis = getCurrentMillis();
            this.cliOptions.outputDir = FilePath(getTempDir()) / "spice" / "output" / toString(millis);
            this.cliOptions.outputPath = this.cliOptions.outputDir / this.cliOptions.mainSourceFile.getFileName();
        } else if this.cliOptions.outputPath.isEmpty() {
            if this.cliOptions.outputPath.isEmpty() {
                this.cliOptions.outputDir = this.cliOptions.outputPath;
                this.cliOptions.outputPath = this.cliOptions.outputDir / this.cliOptions.mainSourceFile.getFileName();
            } else {
                this.cliOptions.outputDir = FilePath(this.cliOptions.outputPath.getParentDir());
            }
        } else {
            this.cliOptions.outputDir = FilePath("./");
            this.cliOptions.outputPath = this.cliOptions.outputDir / this.cliOptions.mainSourceFile.getFileName();
        }

        // Set output file extension
        if this.cliOptions.targetArch == TARGET_WASM32 || this.cliOptions.targetArch == TARGET_WASM64 {
            this.cliOptions.outputPath.replaceExtension("wasm");
        } else if isWindows() {
            this.cliOptions.outputPath.replaceExtension("exe");
        } else {
            this.cliOptions.outputPath.replaceExtension("");
        }

        // Set cache dir
        this.cliOptions.cacheDir = FilePath(getTempDir()) / "spice" / "cache";

        // Create directories in case they not exist yet
        // ToDo
    });*/
}

/**
 * Start the parsing process
 *
 * @param argc Argument count
 * @param argv Argument vector
 * @return Return code
 */
public f<int> Driver.parse(int argc, string[] argv) {
    return this.cliParser.parse(argc, argv);
}

/**
 * Initialize the cli options based on the input of the user
 */
public p Driver.enrich() {
    // Propagate target information
    if this.cliOptions.targetTriple.isEmpty() && this.cliOptions.targetArch.isEmpty() {
        // ToDo: Extend
    }

    // Dump AST, IR and symbol table if all debug output is enabled
    if this.cliOptions.printDebugOutput {
        this.cliOptions.dumpSettings.dumpAST = true;
        this.cliOptions.dumpSettings.dumpIR = true;
        this.cliOptions.dumpSettings.dumpSymbolTable = true;
    }
}

/**
 * Executes the built executable
 */
public p Driver.runBinary() {
    // Print status message
    if this.cliOptions.printDebugOutput {
        print("Running executable ...\n\n");
    }

    // Run executable
    FilePath executablePath = this.cliOptions.outputPath;
    executablePath.makeNative();
    const int exitCode = execCmd(executablePath.toString());
    if exitCode != 0 {
        panic(Error("Your Spice executable exited with non-zero exit code"));
    }
}

/**
 * Add build subcommand to cli interface
 */
p Driver.addBuildSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.addSubcommand("build", "Builds your Spice program and emits an executable");
    subCmd.addAlias("b");

    this.addCompileSubcommandOptions(subCmd);

    // --target-triple
    CliOption<String>& targetOption = subCmd.addOption("--target", this.cliOptions.targetTriple, "Target triple for the emitted executable (for cross-compiling)");
    targetOption.addAlias("--target-triple");
    targetOption.addAlias("-t");
    // --target-arch
    CliOption<String>& targetArchOption = subCmd.addOption("--target-arch", this.cliOptions.targetArch, "Target arch for emitted executable (for cross-compiling)");
    // --target-vendor
    CliOption<String>& targetVendorOption = subCmd.addOption("--target-vendor", this.cliOptions.targetVendor, "Target vendor for emitted executable (for cross-compiling)");
    // --target-os
    CliOption<String>& targetOsOption = subCmd.addOption("--target-os", this.cliOptions.targetOs, "Target OS for emitted executable (for cross-compiling)");

    // --output
    CliOption<FilePath>& outputOption = subCmd.addOption("--output", this.cliOptions.outputPath, "Set the output file path");
    outputOption.addAlias("-o");
    // --debug-info
    CliOption<bool>& debugInfoOption = subCmd.addFlag("--debug-info", this.cliOptions.generateDebugInfo, "Generate debug info");
    debugInfoOption.addAlias("-g");
    // --disable-verifier
    subCmd.addFlag("--disable-verifier", this.cliOptions.disableVerifier, "Disable LLVM module and function verification");
}

/**
 * Add run subcommand to cli interface
 */
p Driver.addRunSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.addSubcommand("run", "Builds your Spice program and runs it immediately");
    subCmd.addAlias("r");

    this.addCompileSubcommandOptions(subCmd);

    // --output
    CliOption<FilePath>& outputOption = subCmd.addOption("--output", this.cliOptions.outputPath, "Set the output file path");
    outputOption.addAlias("-o");
    // --debug-info
    CliOption<bool>& debugInfoOption = subCmd.addFlag("--debug-info", this.cliOptions.generateDebugInfo, "Generate debug info");
    debugInfoOption.addAlias("-g");
    // --disable-verifier
    subCmd.addFlag("--disable-verifier", this.cliOptions.disableVerifier, "Disable LLVM module and function verification");
}

/**
 * Add test subcommand to cli interface
 */
p Driver.addTestSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.addSubcommand("test", "Builds your Spice program and runs all enclosed tests");
    subCmd.addAlias("t");

    this.addCompileSubcommandOptions(subCmd);

    // --debug-info
    CliOption<bool>& debugInfoOption = subCmd.addFlag("--debug-info", this.cliOptions.generateDebugInfo, "Generate debug info");
    debugInfoOption.addAlias("-g");
    // --disable-verifier
    subCmd.addFlag("--disable-verifier", this.cliOptions.disableVerifier, "Disable LLVM module and function verification");
}

/**
 * Add install subcommand to cli interface
 */
p Driver.addInstallSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.addSubcommand("install", "Builds your Spice program and installs it to a directory in the PATH variable");
    subCmd.addAlias("i");

    this.addCompileSubcommandOptions(subCmd);
}

/**
 * Add uninstall subcommand to cli interface
 */
p Driver.addUninstallSubcommand() {
    // Create sub-command itself
    CliSubcommand& subCmd = this.cliParser.addSubcommand("uninstall", "Builds your Spice program and runs it immediately");
    subCmd.addAlias("u");

    this.addCompileSubcommandOptions(subCmd);
}

p Driver.addCompileSubcommandOptions(CliSubcommand& subCmd) {
    const p(string&) buildModeCallback = p(string& buildMode) {
        if buildMode == BUILD_MODE_DEBUG {
            this.cliOptions.buildMode = BuildMode::DEBUG;
        } else if buildMode == BUILD_MODE_RELEASE {
            this.cliOptions.buildMode = BuildMode::RELEASE;
        } else if buildMode == BUILD_MODE_TEST {
            this.cliOptions.buildMode = BuildMode::TEST;
        } else {
            panic(Error("Invalid build mode"));
        }
    };

    // --build-mode
    CliOption<string>& buildModeOption = subCmd.addOption("--build-mode", buildModeCallback, "Build mode (debug, release, test)");
    buildModeOption.addAlias("-m");
    // --llvm-args
    CliOption<String>& llvmArgsOption = subCmd.addOption("--llvm-args", this.cliOptions.llvmArgs, "Additional arguments for LLVM");
    llvmArgsOption.addAlias("-llvm");
    // --jobs
    CliOption<int>& jobsOption = subCmd.addOption("--jobs", this.cliOptions.compileJobCount, "Compile jobs (threads), used for compilation");
    jobsOption.addAlias("-j");
    // --ignore-cache
    subCmd.addFlag("--ignore-cache", this.cliOptions.ignoreCache, "Force re-compilation of all source files");
    // --use-lifetime-markers
    subCmd.addFlag("--use-lifetime-markers", this.cliOptions.useLifetimeMarkers, "Generate lifetime markers to enhance optimizations");

    // Opt levels
    subCmd.addOption("-O0", p(string& _v) { this.cliOptions.optLevel = OptLevel::O0; }, "Disable optimization for the output executable.");
    subCmd.addOption("-O1", p(string& _v) { this.cliOptions.optLevel = OptLevel::O1; }, "Optimization level 1. Only basic optimization is executed.");
    subCmd.addOption("-O2", p(string& _v) { this.cliOptions.optLevel = OptLevel::O2; }, "Optimization level 2. More advanced optimization is applied.");
    subCmd.addOption("-O3", p(string& _v) { this.cliOptions.optLevel = OptLevel::O3; }, "Optimization level 3. Aggressive optimization for best performance.");
    subCmd.addOption("-Os", p(string& _v) { this.cliOptions.optLevel = OptLevel::Os; }, "Optimization level s. Size optimization for output executable.");
    subCmd.addOption("-Oz", p(string& _v) { this.cliOptions.optLevel = OptLevel::Oz; }, "Optimization level z. Aggressive optimization for best size.");
    subCmd.addFlag("-lto", this.cliOptions.useLTO, "Enable link time optimization (LTO)");

    // --debug-output
    CliOption<bool>& debugOutputFlag = subCmd.addFlag("--debug-output", this.cliOptions.printDebugOutput, "Enable debug output");
    debugOutputFlag.addAlias("-d");
    // --dump-cst
    CliOption<bool>& dumpCstFlag = subCmd.addFlag("--dump-cst", this.cliOptions.dumpSettings.dumpCST, "Dump CSTs as serialized string and SVG image");
    dumpCstFlag.addAlias("-cst");
    // --dump-ast
    CliOption<bool>& dumpAstFlag = subCmd.addFlag("--dump-ast", this.cliOptions.dumpSettings.dumpAST, "Dump ASTs as serialized string and SVG image");
    dumpAstFlag.addAlias("-ast");
    // --dump-symtab
    CliOption<bool>& dumpSymtabFlag = subCmd.addFlag("--dump-symtab", this.cliOptions.dumpSettings.dumpSymbolTable, "Dump serialized symbol tables");
    dumpSymtabFlag.addAlias("-symtab");
    // --dump-types
    CliOption<bool>& dumpTypesFlag = subCmd.addFlag("--dump-types", this.cliOptions.dumpSettings.dumpTypes, "Dump all used types");
    dumpTypesFlag.addAlias("-types");
    // --dump-ir
    CliOption<bool>& dumpIrFlag = subCmd.addFlag("--dump-ir", this.cliOptions.dumpSettings.dumpIR, "Dump LLVM-IR");
    dumpIrFlag.addAlias("-ir");
    // --dump-assembly
    CliOption<bool>& dumpAsmFlag = subCmd.addFlag("--dump-assembly", this.cliOptions.dumpSettings.dumpAssembly, "Dump Assembly code");
    dumpAsmFlag.addAlias("-asm");
    dumpAsmFlag.addAlias("-s");
    // --dump-object-file
    CliOption<bool>& dumpObjFlag = subCmd.addFlag("--dump-object-file", this.cliOptions.dumpSettings.dumpObjectFile, "Dump object file");
    dumpObjFlag.addAlias("-obj");

    CliOption<FilePath>& fileOption = subCmd.addOption("<main-source-file>", this.cliOptions.mainSourceFile, "Main source file");
    //fileOption.setRequired();
    //fileOption.check(CliOption::EXISTING_FILE);
}
