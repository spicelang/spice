f<int> main() {
    String test = String("String to be trimmed ");
    printf("'%s'\n", test);
    String trimmed = test.trim();
    printf("'%s'\n", trimmed);
}