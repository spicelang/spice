ext<byte*> malloc(long);
ext free(byte*);

f<int> main() {
    byte* address = malloc(1l);
    *address = (byte) 12;
    free(address);
}