f<int> foo() {
    heap int* ptr = sNew<int>();
    *ptr = 5;
    heap int* ptr2 = ptr;
    return ptr;
}