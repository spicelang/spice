f<int> main() {
    int i = 1;
    i += 2s;
    i *= 2s;
    i /= 2s;
    i -= 2s;
    printf("Result 1: %d\n", i);
    /*i += 223372036854775807l;
    i /= 2l;
    i *= 2l;
    i -= 223372036854775807l;
    printf("Result 2: %d\n", i);*/
}