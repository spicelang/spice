type T int|double;

public type Vector<T> struct {
    public T data
}

public p Vector.setData(T data) {
    this.data = data;
}