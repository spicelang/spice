// Link external functions
ext f<heap byte*> malloc(long);
ext p free(heap byte*);

// Add generic type definitions
type T dyn;

// Enums
type NodeColor enum { RED, BLACK }

/**
 * Node of a Red-Black Tree
 */
type Node<T> struct {
    T data
    heap Node<T>* parent
    heap Node<T>* childLeft
    heap Node<T>* childRight
    NodeColor color
}

inline f<bool> Node.isRoot() {
    return this.parent == nil<heap Node<T>*>;
}

p Node.dump(unsigned int indent = 0) {
    // Dump right child
    if this.childRight != nil<heap Node<T>*> { this.childRight.dump(indent + 4); }
    // Dump node itself
    printf("%s%d %s", String(' ') * indent, this.data, this.color == NodeColor::RED ? "R" : "B");
    // Dump left child
    if this.childLeft != nil<heap Node<T>*> { this.childLeft.dump(indent + 4); }
}

f<heap Node<T>*> createNode<T>(T data) {
    Result<heap Node<T>*> allocResult = sAlloc(sizeof(type Node<T>));
    heap Node<T>* newNode = allocResult.unwrap();
    newNode.data = data;
    newNode.childLeft = nil<heap Node<T>*>;
    newNode.childRight = nil<heap Node<T>*>;
    newNode.color = NodeColor::RED;
    return newNode;
}

/**
 * A Red-Black Tree is a self-balancing search tree, which is used e.g. in the implementation of maps.
 *
 * Insertion time: O(log n)
 * Lookup time: O(log n)
 * Deletion time: O(log n)
 */
public type RedBlackTree<T> struct {
    heap Node<T>* rootNode
}

public p RedBlackTree.ctor() {
    this.rootNode = nil<heap Node<T>*>;
}

public p RedBlackTree.insert(T newItem) {
    heap Node<T>* newNode = createNode<T>(newItem);

}

public p RedBlackTree.insertFixup(heap Node<T>* node) {

}

public p RedBlackTree.dump() {
    if this.rootNode != nil<heap Node<T>*> { this.rootNode.dump(); }
}