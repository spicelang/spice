import "std/iterators/ranges";

f<int> main() {
    //NumberIterator<int> it = range(1, 5);
    for (
        dyn it = range(1l, 10l);
        it.hasNext();
        it.next()
    ) {
        printf("%d\n", it.get());
    }

    /*foreach int i : range(1, 3) {
        printf("%d\n", i);
    }*/
}