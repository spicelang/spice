f<int> main() {
    const dyn variable = 4.3;
    variable = 3.2;
    return 0;
}