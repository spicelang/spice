/**
 * Check if a long is a power of two
 *
 * @param input Input number
 * @return Is power of two
 */
public f<bool> isPowerOfTwo(long input) {
    return (input & (input - 1l)) == 0l;
}