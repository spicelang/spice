// TEST: --output-container=dylib

f<int> add(int a, int b) {
    return a + b;
}