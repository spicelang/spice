import "source1" as s1;

f<int> main() {
    dyn v = s1.Vector<int>{};
    v.setData<int>(12);
    printf("Data: %d\n", v.data);
    v.setData<double>(1.5);
    printf("Data: %d\n", v.data);
}