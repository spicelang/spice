import "std/os/os";
import "std/io/file";

const char PATH_SEPARATOR_UNIX = '/';
const char PATH_SEPARATOR_WINDOWS = '\\';

/**
 * Represents a path to a file or directory on the local file system
 */
public type FilePath struct {
    String path
}

public p FilePath.ctor() {
    this.path = String();
}

public p FilePath.ctor(string pathStr) {
    this.path = String(pathStr);
}

public p FilePath.ctor(const String& pathStr) {
    this.path = pathStr;
}

public p FilePath.ctor(const FilePath& other) {
    this.path = other.path;
}

/**
 * Returns the content of the filepath without modifying.
 *
 * @return The content of the filepath
 */
public f<string> FilePath.toString() {
    return this.path.getRaw();
}

/**
  * Returns the content of the filepath using the given path separator.
  *
  * @param separator The path separator to use
  * @return The content of the filepath using the given path separator
  */
public f<string> FilePath.toStringWithCustomSeparator(char separator) {
    if separator != PATH_SEPARATOR_UNIX {
        this.path.replaceAll(PATH_SEPARATOR_UNIX, separator);
    }
    if separator != PATH_SEPARATOR_WINDOWS {
        this.path.replaceAll(PATH_SEPARATOR_WINDOWS, separator);
    }
    return this.path.getRaw();
}

/**
 * Returns the content of the filepath using the UNIX path separator.
 *
 * @return The content of the filepath using the UNIX path separator
 */
public f<string> FilePath.toGenericString() {
    return this.toStringWithCustomSeparator(PATH_SEPARATOR_UNIX);
}

/**
 * Returns the content of the filepath using the native path separator.
 *
 * @return The content of the filepath using the native path separator
 */
public f<string> FilePath.toNativeString() {
    return this.toStringWithCustomSeparator(isWindows() ? PATH_SEPARATOR_WINDOWS : PATH_SEPARATOR_UNIX);
}

public f<bool> operator==(const FilePath& lhs, const FilePath& rhs) {
    return lhs.path == rhs.path;
}

public f<bool> operator!=(const FilePath& lhs, const FilePath& rhs) {
    return lhs.path != rhs.path;
}

public p operator/=(FilePath& lhs, string rhs) {
    if lhs.path.isEmpty() || rhs[len(rhs) - 1] == PATH_SEPARATOR {
        lhs.path += rhs;
    } else {
        lhs.path += PATH_SEPARATOR;
        lhs.path += rhs;
    }
}

public p operator/=(FilePath& lhs, const String& rhs) {
    lhs /= rhs.getRaw();
}

public p operator/=(FilePath& lhs, const FilePath& rhs) {
    lhs /= rhs.path.getRaw();
}

public f<FilePath> operator/(const FilePath& lhs, string rhs) {
    result = FilePath(lhs);
    result /= rhs;
}

public f<FilePath> operator/(const FilePath& lhs, const String& rhs) {
    result = FilePath(lhs);
    result /= rhs.getRaw();
}

public f<FilePath> operator/(const FilePath& lhs, const FilePath& rhs) {
    result = FilePath(lhs);
    result /= rhs.path.getRaw();
}

/**
 * Checks if the file or directory exists.
 *
 * @return True if the file or directory exists, false otherwise
 */
public f<bool> FilePath.exists() {
    return fileExists(this.path.getRaw());
}