/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "socket" as socket;

f<int> main() {
    socket.Socket s = socket.openServerSocket(8080s);
}*/

// Inspired by: https://www.geeksforgeeks.org/program-for-conways-game-of-life

/*import "std/math/rand" as rand;

const int row = 5;
const int col = 4;

p rowLine() {
    printf("\n");
    for int i = 0; i < col; i++ { printf(" -----"); }
    printf("\n");
}

f<int> countLiveNeighbourCell(int[5][4] a, int r, int c) {
    int count = 0;
    for int i = r - 1; i <= r + 1; i++ {
        for int j = c - 1; j <= c + 1; j++ {
            if (i == r && j == c) || (i < 0 || j < 0) || (i >= row || j >= col) {
                continue;
            }
            if a[i][j] == 1 {
                count++;
            }
        }
    }
    return count;
}

f<int> main() {
    int[5][4] a;
    int[5][4] b;

    // Generate matrix canvas with random values (live and dead cells)
    for int i = 0; i < row; i++ {
        for int j = 0; j < col; j++ {
            a[i][j] = rand.randInt(0, 1);
        }
    }

    printf("Initial state:\n");
    rowLine();
    for int i = 0; i < row; i++ {
        printf(":");
        for int j = 0; j < col; j++ {
            printf("  %d  :", a[i][j]);
        }
        rowLine();
    }
}*/

f<int> main() {
    int i = 0;
    int r = 0;
    int j = 0;
    int c = 0;
    int row = 0;
    int col = 0;
    while(true) {
        if (i == r && j == c) || (i < 0 || j < 0) || (i >= row || j >= col) {
            continue;
        }
        break;
    }
}