// Std imports
import "std/data/vector";

// Own imports
import "bootstrap/util/common-util";
import "bootstrap/ast/ast-nodes";
import "bootstrap/symboltablebuilder/type-chain";
import "bootstrap/symboltablebuilder/qual-type";
import "bootstrap/symboltablebuilder/type-intf";
import "bootstrap/symboltablebuilder/scope-intf";

public type Type struct : IType {
    Vector<TypeChainElement> typeChain
    bool isBaseTypeSigned
}

p Type.ctor(SuperType superType) {
    this.typeChain.pushBack(TypeChainElement(superType));
}

p Type.ctor(SuperType superType, const String& subType) {
    this.typeChain.pushBack(TypeChainElement(superType, subType));
}

p Type.ctor(SuperType superType, const String& subType, unsigned long typeId, const TypeChainElementData& data, const QualTypeList& templateTypes) {
    this.typeChain.pushBack(TypeChainElement(superType, subType, typeId, data, templateTypes));
}

p Type.ctor(TypeChain typeChain) {
    this.typeChain = typeChain.typeChain;
}

/**
 * Get the super type of the current type
 *
 * @return Super type
 */
public f<SuperType> Type.getSuperType() {
    assert !this.typeChain.isEmpty();
    return this.typeChain.back().superType;
}

/**
 * Get the sub type of the current type
 *
 * @return Sub type
 */
public f<const String&> Type.getSubType() {
    assert !this.typeChain.isEmpty();
    const dyn options = [SuperType::TY_STRUCT, SuperType::TY_INTERFACE, SuperType::TY_ENUM, SuperType::TY_GENERIC];
    assert this.isOneOf(options, len(options));
    return this.typeChain.back().subType;
}

/**
 * Get the array size of the current type
 *
 * @return Array size
 */
public f<unsigned int> Type.getArraySize() {
    assert this.isArray();
    return this.typeChain.back().data.arraySize;
}

/**
 * Get the body scope of the current type
 *
 * @return Body scope
 */
public f<IScope*> Type.getBodyScope() {
    const dyn options = [SuperType::TY_STRUCT, SuperType::TY_INTERFACE, SuperType::TY_ENUM, SuperType::TY_GENERIC];
    assert this.isOneOf(options, len(options));
    return this.typeChain.back().data.bodyScope;
}

/**
 * Get the pointer type of the current type as a new type
 *
 * @param node AST node for error messages
 * @return Pointer type of the current type
 */
public f<const Type*> Type.toPtr(const ASTNode* node) {
    if this.is(SuperType::TY_DYN) { panic(Error("Just use the dyn type without '*' instead")); }
    if this.isRef() { panic(Error("Pointers to references are not allowd. Use pointer instead")); }

    // Create new type chain
    TypeChain newTypeChain = this.typeChain;
    newTypeChain.pushBack(TypeChainElement(SuperType::TY_PTR));

    // Register new type or return if already registered
    // ToDo
    return nil<const Type*>;
}

/**
 * Get the reference type of the current type as a new type
 *
 * @param node AST node for error messages
 * @return Reference type of the current type
 */
public f<const Type*> Type.toRef(const ASTNode* node) {
    if this.is(SuperType::TY_DYN) { panic(Error("Just use the dyn type without '&' instead")); }
    if this.isRef() { panic(Error("References to references are not allowd")); }

    // Create new type chain
    TypeChain newTypeChain = this.typeChain;
    newTypeChain.pushBack(TypeChainElement(SuperType::TY_REF));

    // Register new type or return if already registered
    // ToDo
    return nil<const Type*>;
}

/**
 * Get the array type of the current type as a new type
 *
 * @param node AST node for error messages
 * @param size Size of the array
 * @param skipDynCheck Skip check if array base type is dyn
 * @return Array type of the current type
 */
public f<const Type*> Type.toArr(const ASTNode* node, unsigned int size, bool skipDynCheck = false) {
    // Do not allow arrays of dyn
    if !skipDynCheck && this.typeChain.back().superType == SuperType::TY_DYN {
        panic(Error("Just use the dyn type without '[]' instead"));
    }

    // Create new type chain
    TypeChain newTypeChain = this.typeChain;
    TypeChainElementData data = TypeChainElementData{/*arraySize=*/ size, /*bodyScope=*/ nil<IScope*>, /*hasCaptures*/ false};
    newTypeChain.pushBack(TypeChainElement(SuperType::TY_ARRAY, data));

    // Register new type or return if already registered
    // ToDo
    return nil<const Type*>;
}

/**
 * Retrieve the base type of an array or a pointer
 *
 * @return Base type
 */
public f<const Type*> Type.getContained() {
    if this.is(SuperType::TY_STRING) {
        // ToDo
    }

    // Create new type chain
    TypeChain newTypeChain = this.typeChain;
    assert newTypeChain.getSize() > 1;
    newTypeChain.popBack();

    // Register new type or return if already registered
    // ToDo
    return nil<const Type*>;
}

/**
 * Replace the base type with another one
 *
 * @param newBaseType New base type
 * @return The new type
 */
public f<const Type*> Type.replaceBase(const Type* newBaseType) {
    assert !this.typeChain.isEmpty();

    // Create new type
    TypeChain newTypeChain = newBaseType.typeChain;
    const bool doubleRef = newTypeChain.back().superType == SuperType::TY_REF && this.typeChain.back().superType == SuperType::TY_REF;
    foreach unsigned long i = 1ul, const TypeChainElement& element : this.typeChain {
        if !doubleRef || i > 1ul {
            newTypeChain.pushBack(element);
        }
    }

    // Register new type or return if already registered
    // ToDo
    return nil<const Type*>;
}

/**
 * Remove reference wrapper from the current type
 *
 * @return Type without reference wrapper
 */
public f<const Type*> Type.removeReferenceWrapper() {
    return this.isRef() ? this.getContained() : this;
}

/**
 * Return the LLVM type for this symbol type
 *
 * @param sourceFile Referenced source file
 * @return Corresponding LLVM type
 */
public f<llvm::Type> Type.toLLVMType(SourceFile* sourceFile) {
    assert !this.typeChain.isEmpty() && !this.is(SuperType::TY_INVALID);
    llvm::LLVMContext& context = sourceFile.llvmModule.getContext();
}
