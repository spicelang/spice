import "std/type/int";

f<int> main() {
    // toDouble()
    double asDouble = toDouble(123);
    assert asDouble == 123.0;

    // toShort()
    short asShort = toShort(-345);
    assert asShort == -345s;

    // toLong()
    long asLong = toLong(459873);
    assert asLong == 459873l;

    // toByte()
    byte asByte = toByte(12);
    assert asByte == (byte) 12;

    // toChar()
    char asChar = toChar(66);
    assert asChar == 'B';

    // toString()
    String asString = toString(12345);
    assert asString.getRaw() == "12345";

    // toBool()
    bool asBool1 = toBool(1);
    assert asBool1 == true;
    bool asBool2 = toBool(0);
    assert asBool2 == false;

    // isPowerOfTwo()
    assert isPowerOfTwo(16);
    assert !isPowerOfTwo(31);

    printf("All assertions succeeded");
}