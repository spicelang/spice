import "std/iterator/iterable";

// Generic type definitions
type I dyn;
type Numeric int|long|short;

/**
 * A ArrayIterator in Spice can be used to iterate over an arbitrary array
 */
public type ArrayIterator<I> struct : Iterable<I> {
    I* array
    unsigned long size
    unsigned long cursor
}

public p ArrayIterator.ctor(I[] array, unsigned long size) {
    this.array = array;
    this.size = size;
    this.cursor = 0l;
}

/**
 * Returns the current item of the array
 *
 * @return Reference to the current item
 */
public inline f<I&> ArrayIterator.get() {
    unsafe {
        return this.array[this.cursor];
    }
}

public inline f<Pair<unsigned long, I&>> ArrayIterator.getIdx() {
    unsafe {
        return Pair<unsigned long, I&>(this.cursor, this.array[this.cursor]);
    }
}

/**
 * Check if the iterator is valid
 *
 * @return true or false
 */
public inline const f<bool> ArrayIterator.isValid() {
    return this.cursor < this.size;
}

/**
 * Returns the current item of the array and moves the cursor to the next one
 */
public inline p ArrayIterator.next() {
    assert this.isValid();
    this.cursor++;
}

/**
 * Advances the cursor by one
 *
 * @param it ArrayIterator
 */
/*public inline p operator++<I>(ArrayIterator<I>& it) {
    assert it.cursor < it.size- 1;
    it.cursor++;
}*/

/**
 * Move the cursor back by one
 *
 * @param it ArrayIterator
 */
/*public inline p operator--<I>(ArrayIterator<I>& it) {
    assert it.cursor > 0;
    it.cursor--;
}*/

/**
 * Advances the cursor by the given offset
 *
 * @param it ArrayIterator
 * @param offset Offset
 */
/*public inline p operator+=<I, Numeric>(ArrayIterator<I>& it, Numeric offset) {
    assert it.cursor + offset < it.size;
    assert it.cursor + offset >= 0;
    it.cursor += offset;
}*/

/**
 * Move the cursor back by the given offset
 *
 * @param it ArrayIterator
 * @param offset Offset
 */
/*public inline p operator-=<I, Numeric>(ArrayIterator<I>& it, Numeric offset) {
    assert it.cursor - offset < it.size;
    assert it.cursor - offset >= 0;
    it.cursor -= offset;
}*/