f<int> main() {
    dyn[] test = [ "This", "is", "a", "Test" ];
}