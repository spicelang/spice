type Visitor struct {}

type SymbolTable struct {}

type Visitable interface {
    f<bool> accept(Visitor*);
}

type AstNode struct : Visitable {}

type AstEntryNode struct : Visitable {
    AstNode astNode
    SymbolTable* extFunctionScope
    bool takesArgs
}

f<int> main() {
    AstEntryNode entryNode;
    printf("%d", entryNode.takesArgs);
}

/*import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

type ASTNode struct {
    int value
}

p ASTNode.dtor() {
    printf("Dtor called!");
}

f<int> main() {
    DefaultMemoryManager defaultMemoryManager;
    IMemoryManager* memoryManager = &defaultMemoryManager;
    memoryManager.allocate(10l);
    //BlockAllocator<ASTNode> allocator = BlockAllocator<ASTNode>(memoryManager, 10l);
}*/