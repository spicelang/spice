// Constants
public const int TIMEZONE_UTC = 0;

// Structs
type TimeVal struct {
    unsigned long tvSec
    unsigned long tvUsec
}
type TimeZone struct {
    int tzMinutewest
    int tzDsttime
}

// Link external functions
ext f<int> gettimeofday(TimeVal*, TimeZone*);

/**
 * Retrieve seconds since epoch
 */
public f<long> getCurrentSecs() {
    TimeVal time = TimeVal{};
    gettimeofday(&time, nil<TimeZone*>);
    return time.tvSec * 1000l;
}

/**
 * Retrieve milliseconds since epoch
 */
public f<long> getCurrentMillis() {
    TimeVal time = TimeVal{};
    gettimeofday(&time, nil<TimeZone*>);
    return time.tvSec * 1000l + time.tvUsec / 1000l;
}

/**
 * Retrieve microseconds since epoch
 */
public f<long> getCurrentMicros() {
    TimeVal time = TimeVal{};
    gettimeofday(&time, nil<TimeZone*>);
    return 1000000l * time.tvSec + time.tvUsec;
}

/**
 * Check whether a given year is a leap year (Gregorian calendar)
 */
public f<bool> isLeapYear(int year) {
    if year % 400 == 0 {
        return true;
    }
    if year % 100 == 0 {
        return false;
    }
    return year % 4 == 0;
}

/**
 * Return the current UTC year in a fully cross-platform way
 */
public f<int> getCurrentYear() {
    // Seconds since Unix epoch (1970-01-01T00:00:00Z)
    TimeVal time = TimeVal{};
    gettimeofday(&time, nil<TimeZone*>);

    long seconds = time.tvSec;
    long days = seconds / 86400l;

    int year = 1970;

    // Subtract full years until remaining days fit into the current year
    while true {
        const int daysInYear = isLeapYear(year) ? 366 : 365;
        if (days < daysInYear) {
            break;
        }
        days -= daysInYear;
        year++;
    }

    return year;
}
