f<int> main() {
    int i = 1;
    printf("%d", i);
}