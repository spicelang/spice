// TEST: --sanitizer=memory --build-mode=release -g

f<int> main() {
    int i;
    i++;
    printf("%d", i);
}