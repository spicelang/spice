import "std/io/file" as file;

f<int> main() {
    file.File openFile = file.openFile("./test.txt", file.MODE_WRITE);
    openFile.writeChar('A');
    openFile.close();
}