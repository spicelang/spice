import "../exception/ErrorManager";
import "../global/RuntimeModuleManager";
import "../linker/ExternalLinkerInterface";
import "../util/CodeLoc";
import "../util/Timer";
import "../CliInterface";

// Constants
public const string MAIN_FILE_NAME = "root";
public const string LTO_FILE_NAME = "lto-module";

/**
 * The GlobalResourceManager is instantiated at startup of the compiler and serves as distribution point for globally used assets.
 * Other components of the compiler can request the required global resources from the GlobalResourceManager.
 */
public type GlobalResourceManager struct {
    UnorderedMap<String, SourceFile*> sourceFiles
    Vector<ASTNode> astNodes
    const CliOptions& cliOptions
    ExternalLinkerInterface linker
    CacheManager cacheManager
    RuntimeModuleManager runtimeModuleManager
    llvm::Context context
    llvm::IRBuilder builder
    llvm::Module* ltoModule
    llvm::TargetMachine* targetMachine
    Timer totalTimer
    ErrorManager errorManager
}

public p GlobalResourceManager.ctor(const CliOptions& cliOptions) {
    this.cliOptions = cliOptions;
    // ToDo: extend
}

public p GlobalResourceManager.dtor() {
    // Delete all source files
    foreach (const Pair<string, SourceFile *>& sourceFile : sourceFiles) {
        //delete sourceFile.second;
    }

    // Delete target machine
    //delete targetMachine;
}

public f<SourceFile*> GlobalResourceManager.createSourceFile(SourceFile* parent, const String& dependencyName, const FilePath& path, bool isStdFile) {
    // Check if the source file was already added (e.g. by another source file that imports it)
    const String filePathStr = path.toString();
    if sourceFiles.contains(filePathStr) {
        return sourceFiles.get[filePathStr];
    }

    // Create the new source file
    SourceFile* newSourceFile = new SourceFile(parent, dependencyName, path, isStdFile);
    newSourceFile.insert(filePathStr, newSourceFile);
    return newSourceFile;
}