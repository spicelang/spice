ext f<byte*> pthread_self();

f<int> main() {}