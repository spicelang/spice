import "std/io/cli-parser";

type CliOptions struct {
    bool sayHi = false
}

p callback(bool& value) {
    printf("Callback called with value %d\n", value);
}

f<int> main(int argc, string[] argv) {
    CliParser parser = CliParser("Test Program", "This is a simple test program");
    parser.setVersion("v0.1.0");
    parser.setFooter("Copyright (c) Marc Auberer 2021-2023");

    CliOptions options;
    parser.addFlag("--hi", options.sayHi, "Say hi to the user");
    parser.addFlag("--callback", callback, "Call a callback function");
    parser.addFlag("-cb", p(bool& value) {
        printf("CB called with value %d\n", value);
    }, "Call a callback function");

    parser.parse(argc, argv);

    // Print hi if requested
    if options.sayHi {
        printf("Hi!\n");
    }
}