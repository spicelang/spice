type NestedStruct struct {
    double* test
}

type TestStruct struct {
    double f1
    NestedStruct*[3] f2
}

f<int> main() {
    dyn test = 1.24;
    dyn ns = NestedStruct{ &test };
    dyn s = TestStruct{ 5.4, {&ns, &ns, &ns} };
    printf("Double: %f\n", *s.f2[1].test);
}