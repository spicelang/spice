import "std/runtime/iterator_rt";

f<int> main() {
    // Create test array to iterate over
    int[5] a = { 123, 4321, 9876, 321, -99 };

    // Test base functionality
    dyn it = iterate(a, len(a));

    // Test overloaded operators
    it += 3;

    printf("All assertions passed!");
}