import "std/io/cli-subcommand";
import "std/io/cli-option";
import "std/io/filepath";

// Generic types
type T bool|string|String|int|FilePath;
type StrOrConstStrObjRef string|const String&;

public type CliParser struct {
    CliSubcommand rootSubcommand
}

public p CliParser.ctor(string appName, string appDescription = "") {
    this.rootSubcommand = CliSubcommand(nil<CliSubcommand*>, String("v0.1.0"), String(appName), String(appDescription));
}

public p CliParser.ctor(const String& appName, const String& appDescription = String("")) {
    this.rootSubcommand = CliSubcommand(nil<CliSubcommand*>, String("v0.1.0"), appName, appDescription);
}

public p CliParser.setVersion(string versionString) {
    this.rootSubcommand.setVersion(String(versionString));
}

public p CliParser.setVersion(const String& versionString) {
    this.rootSubcommand.setVersion(versionString);
}

public p CliParser.setFooter(string footer) {
    this.rootSubcommand.setFooter(String(footer));
}

public p CliParser.setFooter(const String& footer) {
    this.rootSubcommand.setFooter(footer);
}

public p CliParser.setRootCallback(p() callback) {
    this.rootSubcommand.setCallback(callback);
}

public p CliParser.allowUnknownOptions() {
    this.rootSubcommand.allowUnknownOptions();
}

public f<CliSubcommand&> CliParser.addSubcommand<StrOrConstStrObjRef>(StrOrConstStrObjRef name, StrOrConstStrObjRef description) {
    return this.rootSubcommand.addSubcommand(name, description);
}

#[ignoreUnusedReturnValue]
public f<CliOption<T>&> CliParser.addOption<T, StrOrConstStrObjRef>(StrOrConstStrObjRef name, T& targetVariable, StrOrConstStrObjRef description) {
    return this.rootSubcommand.addOption(name, targetVariable, description);
}

#[ignoreUnusedReturnValue]
public f<CliOption<T>&> CliParser.addOption<T, StrOrConstStrObjRef>(StrOrConstStrObjRef name, p(const T&) callback, StrOrConstStrObjRef description) {
    return this.rootSubcommand.addOption(name, callback, description);
}

#[ignoreUnusedReturnValue]
public f<CliOption<bool>&> CliParser.addFlag<StrOrConstStrObjRef>(StrOrConstStrObjRef name, bool& targetVariable, StrOrConstStrObjRef description) {
   return  this.rootSubcommand.addFlag(name, targetVariable, description);
}

#[ignoreUnusedReturnValue]
public f<CliOption<bool>&> CliParser.addFlag<StrOrConstStrObjRef>(StrOrConstStrObjRef name, p(const bool&) callback, StrOrConstStrObjRef description) {
    return this.rootSubcommand.addFlag(name, callback, description);
}

public f<int> CliParser.parse(unsigned int argc, string[] argv) {
    return this.rootSubcommand.parse(argc, argv);
}