f<int> main() {
    int test = 12;
    test = 13;
    test++;
    printf("%d", test);
}