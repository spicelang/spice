dyn test = true;
dyn invalid;

f<int> main() {
    printf("Bool: %d", test);
}