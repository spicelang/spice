type TLhs dyn;
type TRhs dyn;

// ------------------------------------------ += ------------------------------------------

p plusEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs += rhs;
    assert lhs == expectedResult;
}

p plusEqualTestInnerUnsafe<TRhs>(int* lhs, const TRhs rhs, const int* expectedResult) {
    unsafe {
        lhs += rhs;
    }
    assert lhs == expectedResult;
}

p plusEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    plusEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    plusEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    plusEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    plusEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p plusEqualTest() {
    // Lhs is double
    plusEqualTestOuter<double, double>(1.234, 98.7654, 99.9994, -99.9994, 97.5314, -97.5314);
    // Lhs is int
    plusEqualTestOuter<int, int>(78, 674, 752, -752, 596, -596);
    plusEqualTestOuter<int, short>(78, 7s, 85, -85, -71, 71);
    plusEqualTestOuter<int, long>(78, 2384723l, 2384801, -2384801, 2384645, -2384645);
    // Lhs is short
    plusEqualTestOuter<short, int>(78s, 674, 752s, -752s, 596s, -596s);
    plusEqualTestOuter<short, short>(78s, 7s, 85s, -85s, -71s, 71s);
    plusEqualTestOuter<short, long>(78s, 2384723l, 25505s, -25505s, 25349s, -25349s);
    // Lhs is long
    plusEqualTestOuter<long, int>(78l, 674, 752l, -752l, 596l, -596l);
    plusEqualTestOuter<long, short>(78l, 7s, 85l, -85l, -71l, 71l);
    plusEqualTestOuter<long, long>(78l, 2384723l, 2384801l, -2384801l, 2384645l, -2384645l);
    // Lhs is char
    plusEqualTestInner<char, int>('A', 5, 'F');
    plusEqualTestInner<char, int>('A', -5, '<');
    // Lhs is ptr
    int[5] input = [0, 0, 0, 0, 0];
    plusEqualTestInnerUnsafe(&input[2], 2, &input[4]);
    plusEqualTestInnerUnsafe(&input[2], -2, &input[0]);
    plusEqualTestInnerUnsafe(&input[2], 2s, &input[4]);
    plusEqualTestInnerUnsafe(&input[2], -2s, &input[0]);
    plusEqualTestInnerUnsafe(&input[2], 2l, &input[4]);
    plusEqualTestInnerUnsafe(&input[2], -2l, &input[0]);
}

// ------------------------------------------ -= ------------------------------------------

p minusEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs -= rhs;
    assert lhs == expectedResult;
}

p minusEqualTestInnerUnsafe<TRhs>(int* lhs, const TRhs rhs, const int* expectedResult) {
    unsafe {
        lhs -= rhs;
    }
    assert lhs == expectedResult;
}

p minusEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    minusEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    minusEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    minusEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    minusEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p minusEqualTest() {
    // Lhs is double
    minusEqualTestOuter<double, double>(1.234, 98.7654, -97.5314, 97.5314, -99.9994, 99.9994);
    // Lhs is int
    minusEqualTestOuter<int, int>(78, 674, -596, 596, -752, 752);
    minusEqualTestOuter<int, short>(78, 7s, 71, -71, -85, 85);
    minusEqualTestOuter<int, long>(78, 2384723l, -2384645, 2384645, -2384801, 2384801);
    // Lhs is short
    minusEqualTestOuter<short, int>(78s, 674, -596s, 596s, -752s, 752s);
    minusEqualTestOuter<short, short>(78s, 7s, 71s, -71s, -85s, 85s);
    // Note: wrap-around consistent with short semantics
    minusEqualTestOuter<short, long>(78s, 2384723l, cast<short>(78s - 2384723l), cast<short>(-78s - -2384723l), cast<short>(-78s - 2384723l), cast<short>(78s - -2384723l));
    // Lhs is long
    minusEqualTestOuter<long, int>(78l, 674, -596l, 596l, -752l, 752l);
    minusEqualTestOuter<long, short>(78l, 7s, 71l, -71l, -85l, 85l);
    minusEqualTestOuter<long, long>(78l, 2384723l, -2384645l, 2384645l, -2384801l, 2384801l);
    // Lhs is char
    minusEqualTestInner<char, int>('A', 5, '<');
    minusEqualTestInner<char, int>('A', -5, 'F');
    // Lhs is ptr
    int[5] input = [0, 0, 0, 0, 0];
    minusEqualTestInnerUnsafe(&input[2], 2, &input[0]);
    minusEqualTestInnerUnsafe(&input[2], -2, &input[4]);
    minusEqualTestInnerUnsafe(&input[2], 2s, &input[0]);
    minusEqualTestInnerUnsafe(&input[2], -2s, &input[4]);
    minusEqualTestInnerUnsafe(&input[2], 2l, &input[0]);
    minusEqualTestInnerUnsafe(&input[2], -2l, &input[4]);
}

// ------------------------------------------ *= ------------------------------------------

p mulEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs *= rhs;
    assert lhs == expectedResult;
}

p mulEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    mulEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    mulEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    mulEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    mulEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p mulEqualTest() {
    // Lhs double
    mulEqualTestOuter<double, double>(1.5, 2.0, 3.0, 3.0, -3.0, -3.0);
    // Lhs int
    mulEqualTestOuter<int, int>(6, 7, 42, 42, -42, -42);
    mulEqualTestOuter<int, short>(6, 3s, 18, 18, -18, -18);
    mulEqualTestOuter<int, long>(6, 5l, 30, 30, -30, -30);
    // Lhs short
    mulEqualTestOuter<short, int>(6s, 7, 42s, 42s, -42s, -42s);
    mulEqualTestOuter<short, short>(6s, 3s, 18s, 18s, -18s, -18s);
    // Note: wrap-around consistent with short semantics
    mulEqualTestOuter<short, long>(200s, 2000l, cast<short>(200 * 2000), cast<short>(-200 * -2000), cast<short>(-200 * 2000), cast<short>(200 * -2000));
    // Lhs long
    mulEqualTestOuter<long, int>(6l, 7, 42l, 42l, -42l, -42l);
    mulEqualTestOuter<long, short>(6l, 3s, 18l, 18l, -18l, -18l);
    mulEqualTestOuter<long, long>(6l, 5l, 30l, 30l, -30l, -30l);
}

// ------------------------------------------ /= ------------------------------------------

p divEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs /= rhs;
    assert lhs == expectedResult;
}

p divEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    divEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    divEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    divEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    divEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p divEqualTest() {
    // Lhs double
    divEqualTestOuter<double, double>(9.0, 3.0, 3.0, 3.0, -3.0, -3.0);
    // Lhs int
    divEqualTestOuter<int, int>(42, 7, 6, 6, -6, -6);
    divEqualTestOuter<int, short>(42, 3s, 14, 14, -14, -14);
    divEqualTestOuter<int, long>(42, 6l, 7, 7, -7, -7);
    // Lhs short
    divEqualTestOuter<short, int>(42s, 7, 6s, 6s, -6s, -6s);
    divEqualTestOuter<short, short>(42s, 3s, 14s, 14s, -14s, -14s);
    divEqualTestOuter<short, long>(100s, 25l, 4s, 4s, -4s,- 4s);
    // Lhs long
    divEqualTestOuter<long, int>(42l, 7, 6l, 6l, -6l, -6l);
    divEqualTestOuter<long, short>(42l, 3s, 14l, 14l, -14l, -14l);
    divEqualTestOuter<long, long>(42l, 6l, 7l, 7l, -7l, -7l);
}

// ------------------------------------------ %= ------------------------------------------

p remEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs %= rhs;
    assert lhs == expectedResult;
}

p remEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    remEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    remEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    remEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    remEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p remEqualTest() {
    // Lhs double
    remEqualTestOuter<double, double>(9.0, 3.0, 0.0, 0.0, 0.0, 0.0);
    // Lhs int
    remEqualTestOuter<int, int>(42, 7, -0, -0, 0, 0);
    remEqualTestOuter<int, short>(42, 8s, 2, -2, -2, 2);
    remEqualTestOuter<int, long>(42, 9l, 6, -6, -6, 6);
    // Lhs short
    remEqualTestOuter<short, int>(42s, 7, -0s, -0s, 0s, 0s);
    remEqualTestOuter<short, short>(42s, 8s, 2s, -2s, -2s, 2s);
    remEqualTestOuter<short, long>(100s, 26l, 22s, -22s, -22s, 22s);
    // Lhs long
    remEqualTestOuter<long, int>(42l, 7, -0l, -0l, 0l, 0l);
    remEqualTestOuter<long, short>(42l, 10s, 2l, -2l, -2l, 2l);
    remEqualTestOuter<long, long>(10932847123l, 234324l, 226579l, -226579l, -226579l, 226579l);
    // Lhs byte
    remEqualTestInner<byte, byte>(cast<byte>(42), cast<byte>(41), cast<byte>(1));
}

// ------------------------------------------ <<= -----------------------------------------

p shlEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs <<= rhs;
    assert lhs == expectedResult;
}

p shlEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2) {
    shlEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    shlEqualTestInner(-lhs, rhs, expectedResult2);  // Lhs -, Rhs +
}

p shlEqualTest() {
    // Lhs int
    shlEqualTestOuter<int, int>(5, 3, 40, -40);
    shlEqualTestOuter<int, short>(5, 2s, 20, -20);
    shlEqualTestOuter<int, long>(5, 4l, 80, -80);
    // Lhs short
    shlEqualTestOuter<short, int>(8s, 2, 32s, -32s);
    shlEqualTestOuter<short, short>(8s, 1s, 16s, -16s);
    shlEqualTestOuter<short, long>(8s, 6l, 512s, -512s);
    // Lhs long
    shlEqualTestOuter<long, int>(7l, 7, 896l, -896l);
    shlEqualTestOuter<long, short>(7l, 10s, 7168l, -7168l);
    shlEqualTestOuter<long, long>(1234876l, 21l, 2589722673152l, -2589722673152l);
    // Lhs byte
    shlEqualTestInner<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(84));
}

// ------------------------------------------ >>= -----------------------------------------

p shrEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs >>= rhs;
    assert lhs == expectedResult;
}

p shrEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2) {
    shrEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    shrEqualTestInner(-lhs, rhs, expectedResult2);  // Lhs -, Rhs +
}

p shrEqualTest() {
    // Lhs int
    shrEqualTestOuter<int, int>(5, 3, 0, -1);
    shrEqualTestOuter<int, short>(5, 2s, 1, -2);
    shrEqualTestOuter<int, long>(5, 1l, 2, -3);
    // Lhs short
    shrEqualTestOuter<short, int>(8s, 2, 2s, -2s);
    shrEqualTestOuter<short, short>(8s, 1s, 4s, 32764s);
    shrEqualTestOuter<short, long>(8s, 3l, 1s, -1s);
    // Lhs long
    shrEqualTestOuter<long, int>(23425l, 7, 183l, -184l);
    shrEqualTestOuter<long, short>(34587334534l, 10s, 33776693l, -33776694l);
    shrEqualTestOuter<long, long>(1234876l, 21l, 0l, -1l);
    // Lhs byte
    shrEqualTestInner<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(21));
}

// ------------------------------------------ &= ------------------------------------------

p andEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs &= rhs;
    assert lhs == expectedResult;
}

p andEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    andEqualTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p andEqualTest() {
    // Lhs int
    andEqualTestOuter<int, int>(5, 3, 1);
    andEqualTestOuter<int, short>(5, 2s, 0);
    andEqualTestOuter<int, long>(5, 1l, 1);
    // Lhs short
    andEqualTestOuter<short, int>(8s, 2, 0s);
    andEqualTestOuter<short, short>(8s, 1s, 0s);
    andEqualTestOuter<short, long>(8s, 3l, 0s);
    // Lhs long
    andEqualTestOuter<long, int>(23425l, 7, 1l);
    andEqualTestOuter<long, short>(34587334534l, 10s, 2l);
    andEqualTestOuter<long, long>(1234876l, 21l, 20l);
    // Lhs byte
    andEqualTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(0));
}

// ------------------------------------------ |= ------------------------------------------

p orEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs |= rhs;
    assert lhs == expectedResult;
}

p orEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    orEqualTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p orEqualTest() {
    // Lhs int
    orEqualTestOuter<int, int>(5, 3, 7);
    orEqualTestOuter<int, short>(5, 2s, 7);
    orEqualTestOuter<int, long>(5, 1l, 5);
    // Lhs short
    orEqualTestOuter<short, int>(8s, 2, 10s);
    orEqualTestOuter<short, short>(8s, 1s, 9s);
    orEqualTestOuter<short, long>(8s, 3l, 11s);
    // Lhs long
    orEqualTestOuter<long, int>(23425l, 7, 23431l);
    orEqualTestOuter<long, short>(34587334534l, 10s, 34587334542l);
    orEqualTestOuter<long, long>(1234876l, 21l, 1234877l);
    // Lhs byte
    orEqualTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(43));
}

// ------------------------------------------ ^= ------------------------------------------

p xorEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs ^= rhs;
    assert lhs == expectedResult;
}

p xorEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    xorEqualTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p xorEqualTest() {
    // Lhs int
    xorEqualTestOuter<int, int>(5, 3, 6);
    xorEqualTestOuter<int, short>(5, 2s, 7);
    xorEqualTestOuter<int, long>(5, 1l, 4);
    // Lhs short
    xorEqualTestOuter<short, int>(8s, 2, 10s);
    xorEqualTestOuter<short, short>(8s, 1s, 9s);
    xorEqualTestOuter<short, long>(8s, 3l, 11s);
    // Lhs long
    xorEqualTestOuter<long, int>(23425l, 7, 23430l);
    xorEqualTestOuter<long, short>(34587334534l, 10s, 34587334540l);
    xorEqualTestOuter<long, long>(1234876l, 21l, 1234857l);
    // Lhs byte
    xorEqualTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(43));
}

// ------------------------------------------ ^ ------------------------------------------

p bitwiseXorTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs ^ rhs;
    printf("actualResult: %lld, expectedResult: %lld\n", actualResult, expectedResult);
    assert actualResult == expectedResult;
}

p bitwiseXorTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    bitwiseXorTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p bitwiseXorTest() {
    // Lhs int
    bitwiseXorTestOuter<int, int>(5, 3, 6);
    // Lhs short
    bitwiseXorTestOuter<short, short>(8s, 1s, 9s);
    // Lhs long
    bitwiseXorTestOuter<long, long>(1234876l, 21l, 1234857l);
    // Lhs byte
    bitwiseXorTestOuter<byte, byte>(cast<byte>(15), cast<byte>(23), cast<byte>(24));
    // Lhs bool
    bitwiseXorTestOuter<bool, bool>(false, false, false);
    bitwiseXorTestOuter<bool, bool>(false, true, true);
    bitwiseXorTestOuter<bool, bool>(true, false, true);
    bitwiseXorTestOuter<bool, bool>(true, true, false);
}

// ------------------------------------------ | ------------------------------------------

p bitwiseOrTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs | rhs;
    assert actualResult == expectedResult;
}

p bitwiseOrTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    bitwiseOrTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p bitwiseOrTest() {
    // Lhs int
    bitwiseOrTestOuter<int, int>(5, 3, 7);
    // Lhs short
    bitwiseOrTestOuter<short, short>(8s, 1s, 9s);
    // Lhs long
    bitwiseOrTestOuter<long, long>(1234876l, 21l, 1234877l);
    // Lhs byte
    bitwiseOrTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(43));
    // Lhs bool
    bitwiseOrTestOuter<bool, bool>(false, false, false);
    bitwiseOrTestOuter<bool, bool>(false, true, true);
    bitwiseOrTestOuter<bool, bool>(true, false, true);
    bitwiseOrTestOuter<bool, bool>(true, true, true);
}

// ------------------------------------------ & ------------------------------------------

p bitwiseAndTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs & rhs;
    printf("actualResult: %lld, expectedResult: %lld\n", actualResult, expectedResult);
    assert actualResult == expectedResult;
}

p bitwiseAndTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    bitwiseAndTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p bitwiseAndTest() {
    // Lhs int
    bitwiseAndTestOuter<int, int>(5, 3, 1);
    // Lhs short
    bitwiseAndTestOuter<short, short>(8s, 1s, 0s);
    // Lhs long
    bitwiseAndTestOuter<long, long>(1234876l, 21l, 20l);
    // Lhs byte
    bitwiseAndTestOuter<byte, byte>(cast<byte>(15), cast<byte>(23), cast<byte>(7));
    // Lhs bool
    bitwiseAndTestOuter<bool, bool>(false, false, false);
    bitwiseAndTestOuter<bool, bool>(false, true, false);
    bitwiseAndTestOuter<bool, bool>(true, false, false);
    bitwiseAndTestOuter<bool, bool>(true, true, true);
}

f<int> main() {
    plusEqualTest();  // +=
    minusEqualTest(); // -=
    mulEqualTest();   // *=
    divEqualTest();   // /=
    remEqualTest();   // %=
    shlEqualTest();   // <<=
    shrEqualTest();   // >>=
    andEqualTest();   // &=
    orEqualTest();    // |=
    xorEqualTest();   // ^=
    bitwiseOrTest();  // |
    bitwiseXorTest(); // ^
    bitwiseAndTest(); // &
    // ToDo: Extend

    printf("All assertions passed!");
}