import "std/iterators/ranges";

f<int> main() {
    //dyn it = range(1, 5);
    //assert it.hasNext();
    //assert it.next() == 2;
    foreach int i : range(1, 5) {
        printf("%d\n", i);
    }
}