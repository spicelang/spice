f<int> main() {
    int& ref;
    ref = 123;
}