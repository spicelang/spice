f<int> greatestCommonDivisor(int a, int b) {
    while b != 0 {
        int temp = b;
        b = a % b;
        a = temp;
    }
    return a;
}

f<int> main() {
    int a = 56;
    int b = 98;
    int gcd = greatestCommonDivisor(a, b);
    printf("GCD of %d and %d is %d.", a, b, gcd);
}
