f<string> getTestString(int _arg0, double _arg1, bool _arg2 = false, double _arg3 = 1.34) {
    return "Test";
}

f<int> main() {
    printf("Result: %s\n", getTestString(1, 3.4, true));
}