ext f<unsigned int> snprintf(string, unsigned long, string, ...);

f<int> main() {
    double input = 3.141590;
    char[100] str;
    snprintf(cast<string>(str), sizeof(str), "%f", input);
    printf("%s", str);
}