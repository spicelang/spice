// Std imports
import "std/data/stack";

// Own imports
//import "bootstrap/compiler-pass";
import "bootstrap/lexer/lexer";
import "bootstrap/lexer/token";
import "bootstrap/ast/ast-nodes";
import "bootstrap/util/block-allocator";

// Generic types
type T dyn;

public type Parser struct {
    //compose CompilerPass compilerPass
    Lexer& lexer
    Stack<ASTNode*> parentStack
    BlockAllocator<ASTNode> astNodeAlloc // ToDo: Remove and use allocator from resource manager via compilerPass
}

public p Parser.ctor(Lexer& lexer) {
    this.lexer = lexer;
}

/*public p Parser.ctor(SourceFile* sourceFile, Lexer& lexer) {
    this.lexer = lexer;
}*/

f<T*> Parser.createNode<T>() {
    ASTNode* parent = nil<ASTNode*>;
    const bool isRootNode = this.parentStack.isEmpty();
    if !isRootNode {
        parent = this.parentStack.top();
    }

    // Create the new node
    //T* node = this.resourceManager.astNodeAlloc.allocate(T(this.lexer.getCodeLoc()));
    T* node = this.astNodeAlloc.allocate(T(this.lexer.getCodeLoc()));

    // If this is not the entry node, we need to add the new node to its parent
    if !isRootNode {
        parent.addChild(node);
    }

    // This node is the parent for its children
    this.parentStack.push(node);

    return node;
}

f<T*> Parser.concludeNode<T>(T* node) {
    assert !this.parentStack.isEmpty();
    assert this.parentStack.top() == node;
    this.parentStack.pop();
    return node;
}

inline f<bool> Parser.currentTokenIs(TokenType expectedTokenType) {
    return this.lexer.getToken().tokenType == expectedTokenType;
}

f<bool> Parser.currentTokenIsOneOf(TokenType[] expectedTokenTypeArray, unsigned long size) {
    for unsigned long i = 0l; i < size; i++ {
        if this.currentTokenIs(expectedTokenTypeArray[i]) {
            return true;
        }
    }
    return false;
}

public f<ASTEntryNode*> Parser.parse() {
    dyn entryNode = this.createNode<ASTEntryNode>();

    while !this.currentTokenIs(TokenType::EOF) {
        this.parseStmt();
    }

    return this.concludeNode(entryNode);
}

public f<ASTMainFctDefNode*> Parser.parseMainFctDef() {
    dyn mainFctDefNode = this.createNode<ASTMainFctDefNode>();

    // Parse topLevelDefAttr
    if this.currentTokenIs(TokenType::FCT_ATTR_PREAMBLE) {
        this.parseTopLevelDefAttr();
    }

    // Parse specifierLst
    if !this.currentTokenIs(TokenType::F) {
        this.parseSpecifierLst();
    }

    // Consume expected tokens 'f<int> main'
    this.lexer.expect(TokenType::F);
    this.lexer.expect(TokenType::LESS);
    this.lexer.expect(TokenType::TYPE_INT);
    this.lexer.expect(TokenType::GREATER);
    this.lexer.expect(TokenType::MAIN);

    // Parse praamLst
    this.lexer.expect(TokenType::LPAREN);
    if !this.currentTokenIs(TokenType::RPAREN) {
        this.parseParamLst();
    }
    this.lexer.expect(TokenType::RPAREN);

    // Parse stmtLst
    this.parseStmtLst();

    return this.concludeNode(mainFctDefNode);
}

public f<ASTFctDefNode*> Parser.parseFctDef() {
    dyn fctDefNode = this.createNode<ASTFctDefNode>();

    // Parse topLevelDefAttr
    if this.currentTokenIs(TokenType::FCT_ATTR_PREAMBLE) {
        this.parseTopLevelDefAttr();
    }

    // Parse specifierLst
    if !this.currentTokenIs(TokenType::F) {
        this.parseSpecifierLst();
    }

    this.lexer.expect(TokenType::F);
    this.lexer.expect(TokenType::LESS);
    this.parseDataType();
    this.lexer.expect(TokenType::GREATER);
    this.parseFctName();

    // Parse typeLst (template type list)
    if this.currentTokenIs(TokenType::LESS) {
        this.lexer.expect(TokenType::LESS);
        this.parseTypeLst();
        this.lexer.expect(TokenType::GREATER);
    }

    // Parse paramLst
    this.lexer.expect(TokenType::LPAREN);
    if !this.currentTokenIs(TokenType::RPAREN) {
        this.parseParamLst();
    }
    this.lexer.expect(TokenType::RPAREN);

    // Parse stmtLst
    this.parseStmtLst();

    return this.concludeNode(fctDefNode);
}

public f<ASTProcDefNode*> Parser.parseProcDef() {
    dyn procDefNode = this.createNode<ASTProcDefNode>();

    // Parse topLevelDefAttr
    if this.currentTokenIs(TokenType::FCT_ATTR_PREAMBLE) {
        this.parseTopLevelDefAttr();
    }

    // Parse specifierLst
    if !this.currentTokenIs(TokenType::P) {
        this.parseSpecifierLst();
    }

    this.lexer.expect(TokenType::P);
    this.parseFctName();

    // Parse typeLst (template type list)
    if this.currentTokenIs(TokenType::LESS) {
        this.lexer.expect(TokenType::LESS);
        this.parseTypeLst();
        this.lexer.expect(TokenType::GREATER);
    }

    // Parse paramLst
    this.lexer.expect(TokenType::LPAREN);
    if !this.currentTokenIs(TokenType::RPAREN) {
        this.parseParamLst();
    }
    this.lexer.expect(TokenType::RPAREN);

    // Parse stmtLst
    this.parseStmtLst();

    return this.concludeNode(procDefNode);
}

f<ASTFctNameNode*> Parser.parseFctName() {
    dyn fctNameNode = this.createNode<ASTFctNameNode>();

    if this.currentTokenIs(TokenType::OPERATOR) {
        this.lexer.expect(TokenType::OPERATOR);
        // ToDo: consume overloadable op correctly
        this.lexer.advance();
    } else {
        if this.currentTokenIs(TokenType::TYPE_IDENTIFIER) {
            this.lexer.expect(TokenType::TYPE_IDENTIFIER);
            this.lexer.expect(TokenType::DOT);
        }
        this.lexer.expect(TokenType::IDENTIFIER);
    }

    return this.concludeNode(fctNameNode);
}

f<ASTStructDefNode*> Parser.parseStructDef() {
    dyn structDefNode = this.createNode<ASTStructDefNode>();

    // Parse topLevelDefAttr
    if this.currentTokenIs(TokenType::FCT_ATTR_PREAMBLE) {
        this.parseTopLevelDefAttr();
    }

    // Parse specifierLst
    if !this.currentTokenIs(TokenType::TYPE) {
        this.parseSpecifierLst();
    }

    this.lexer.expect(TokenType::TYPE);
    this.lexer.expect(TokenType::TYPE_IDENTIFIER);

    // Parse typeLst (template type list)
    if this.currentTokenIs(TokenType::LESS) {
        this.lexer.expect(TokenType::LESS);
        this.parseTypeLst();
        this.lexer.expect(TokenType::GREATER);
    }

    this.lexer.expect(TokenType::STRUCT);

    // Parse typeLst (implemented interfaces)
    if this.currentTokenIs(TokenType::COLON) {
        this.lexer.expect(TokenType::COLON);
        this.parseTypeLst();
    }

    // Parse fieldLst
    this.lexer.expect(TokenType::LBRACE);
    while !this.currentTokenIs(TokenType::RBRACE) {
        this.parseField();
    }
    this.lexer.expect(TokenType::RBRACE);

    return this.concludeNode(structDefNode);
}

f<ASTInterfaceDefNode*> Parser.parseInterfaceDef() {
    dyn interfaceDefNode = this.createNode<ASTInterfaceDefNode>();

    // Parse topLevelDefAttr
    if this.currentTokenIs(TokenType::FCT_ATTR_PREAMBLE) {
        this.parseTopLevelDefAttr();
    }

    // Parse specifierLst
    if !this.currentTokenIs(TokenType::TYPE) {
        this.parseSpecifierLst();
    }

    this.lexer.expect(TokenType::TYPE);
    this.lexer.expect(TokenType::TYPE_IDENTIFIER);

    // Parse typeLst (template type list)
    if this.currentTokenIs(TokenType::LESS) {
        this.lexer.expect(TokenType::LESS);
        this.parseTypeLst();
        this.lexer.expect(TokenType::GREATER);
    }

    this.lexer.expect(TokenType::INTERFACE);

    // Parse signatures
    this.lexer.expect(TokenType::LBRACE);
    do {
        this.parseSignature();
    } while !this.currentTokenIs(TokenType::RBRACE);
    this.lexer.expect(TokenType::RBRACE);

    return this.concludeNode(interfaceDefNode);
}

f<ASTEnumDefNode*> Parser.parseEnumDef() {
    dyn enumDefNode = this.createNode<ASTEnumDefNode>();

    // Parse specifierLst
    if !this.currentTokenIs(TokenType::TYPE) {
        this.parseSpecifierLst();
    }

    this.lexer.expect(TokenType::TYPE);
    this.lexer.expect(TokenType::TYPE_IDENTIFIER);
    this.lexer.expect(TokenType::ENUM);

    // Parse enumItemLst
    this.lexer.expect(TokenType::LBRACE);
    this.parseEnumItemLst();
    this.lexer.expect(TokenType::RBRACE);

    return this.concludeNode(enumDefNode);
}

f<ASTGenericTypeDefNode*> Parser.parseGenericTypeDef() {
    dyn genericTypeDefNode = this.createNode<ASTGenericTypeDefNode>();

    this.lexer.expect(TokenType::TYPE);
    this.lexer.expect(TokenType::TYPE_IDENTIFIER);
    this.parseTypeAltsLst();
    this.lexer.expect(TokenType::SEMICOLON);

    return this.concludeNode(genericTypeDefNode);
}

f<ASTAliasDefNode*> Parser.parseAliasDef() {
    dyn aliasDefNode = this.createNode<ASTAliasDefNode>();

    // Parse specifierLst
    if !this.currentTokenIs(TokenType::TYPE) {
        this.parseSpecifierLst();
    }

    this.lexer.expect(TokenType::TYPE);
    this.lexer.expect(TokenType::TYPE_IDENTIFIER);
    this.lexer.expect(TokenType::ALIAS);
    this.parseDataType();
    this.lexer.expect(TokenType::SEMICOLON);

    return this.concludeNode(aliasDefNode);
}

f<ASTGlobalVarDefNode*> Parser.parseGlobalVarDef() {
    dyn globalVarDefNode = this.createNode<ASTGlobalVarDefNode>();

    this.parseDataType();
    this.lexer.expect(TokenType::TYPE_IDENTIFIER);

    // Parse initializer
    if !this.currentTokenIs(TokenType::ASSIGN) {
        this.lexer.expect(TokenType::ASSIGN);
        this.parseConstant();
    }

    this.lexer.expect(TokenType::SEMICOLON);

    return this.concludeNode(globalVarDefNode);
}

f<ASTExtDeclNode*> Parser.parseExtDecl() {
    dyn extDeclNode = this.createNode<ASTExtDeclNode>();

    // Parse topLevelDefAttr
    if this.currentTokenIs(TokenType::FCT_ATTR_PREAMBLE) {
        this.parseTopLevelDefAttr();
    }

    this.lexer.expect(TokenType::EXT);

    // Parse parse function prefix / procedure prefix
    if this.currentTokenIs(TokenType::F) {
        this.lexer.expect(TokenType::F);
        this.lexer.expect(TokenType::LESS);
        this.parseDataType();
        this.lexer.expect(TokenType::GREATER);
    } else {
        this.lexer.expect(TokenType::P);
    }

    // Parse external function name
    if this.currentTokenIs(TokenType::IDENTIFIER) {
        this.lexer.expect(TokenType::IDENTIFIER);
    } else {
        this.lexer.expect(TokenType::TYPE_IDENTIFIER);
    }

    // Parse typeLst (param list)
    this.lexer.expect(TokenType::LPAREN);
    if !this.currentTokenIs(TokenType::RPAREN) {
        this.parseTypeLst();
        if this.currentTokenIs(TokenType::ELLIPSIS) {
            this.lexer.expect(TokenType::ELLIPSIS);
        }
    }
    this.lexer.expect(TokenType::RPAREN);

    this.lexer.expect(TokenType::SEMICOLON);

    return this.concludeNode(extDeclNode);
}

f<ASTImportDefNode*> Parser.parseImportDef() {
    dyn importDefNode = this.createNode<ASTImportDefNode>();

    this.lexer.expect(TokenType::IMPORT);
    this.lexer.expect(TokenType::STRING_LIT);

    if this.currentTokenIs(TokenType::AS) {
        this.lexer.expect(TokenType::AS);
        this.lexer.expect(TokenType::IDENTIFIER);
    }
    this.lexer.expect(TokenType::SEMICOLON);

    return this.concludeNode(importDefNode);
}

f<ASTUnsafeBlockNode*> Parser.parseUnsafeBlock() {
    dyn unsafeBlockNode = this.createNode<ASTUnsafeBlockNode>();

    this.lexer.expect(TokenType::UNSAFE);
    this.parseStmtLst();

    return this.concludeNode(unsafeBlockNode);
}

f<ASTForLoopNode*> Parser.parseForLoop() {
    dyn forLoopNode = this.createNode<ASTForLoopNode>();

    this.lexer.expect(TokenType::FOR);

    // Parse head
    if this.currentTokenIs(TokenType::LPAREN) {
        this.lexer.expect(TokenType::LPAREN);
        this.parseForHead();
        this.lexer.expect(TokenType::RPAREN);
    } else {
        this.parseAssignExpr();
    }

    // Parse stmtLst
    this.parseStmtLst();

    return this.concludeNode(forLoopNode);
}

p Parser.parseForHead() {
    this.parseDeclStmt();
    this.lexer.expect(TokenType::SEMICOLON);
    this.parseAssignExpr();
    this.lexer.expect(TokenType::SEMICOLON);
    this.parseAssignExpr();
}

f<ASTForeachLoopNode*> Parser.parseForeachLoop() {
    dyn foreachLoopNode = this.createNode<ASTForeachLoopNode>();

    this.lexer.expect(TokenType::FOREACH);

    // Parse head
    if this.currentTokenIs(TokenType::LPAREN) {
        this.lexer.expect(TokenType::LPAREN);
        this.parseForeachHead();
        this.lexer.expect(TokenType::RPAREN);
    } else {
        this.parseAssignExpr();
    }

    // Parse stmtLst
    this.lexer.expect(TokenType::LBRACE);
    this.parseStmtLst();
    this.lexer.expect(TokenType::RBRACE);

    return this.concludeNode(foreachLoopNode);
}

p Parser.parseForeachHead() {
    this.parseDeclStmt();
    if this.currentTokenIs(TokenType::COMMA) {
        this.lexer.expect(TokenType::COMMA);
        this.parseDeclStmt();
    }
    this.lexer.expect(TokenType::COLON);
    this.parseAssignExpr();
}

f<ASTWhileLoopNode*> Parser.parseWhileLoop() {
    dyn whileLoopNode = this.createNode<ASTWhileLoopNode>();

    this.lexer.expect(TokenType::WHILE);

    // Parse head
    this.parseAssignExpr();

    // Parse stmtLst
    this.parseStmtLst();

    return this.concludeNode(whileLoopNode);
}

f<ASTDoWhileLoopNode*> Parser.parseDoWhileLoop() {
    dyn doWhileLoopNode = this.createNode<ASTDoWhileLoopNode>();

    this.lexer.expect(TokenType::DO);

    // Parse stmtLst
    this.parseStmtLst();

    // Parse foot
    this.lexer.expect(TokenType::WHILE);
    this.parseAssignExpr();
    this.lexer.expect(TokenType::SEMICOLON);

    return this.concludeNode(doWhileLoopNode);
}

f<ASTIfStmtNode*> Parser.parseIfStmt() {
    dyn ifStmtNode = this.createNode<ASTIfStmtNode>();

    this.lexer.expect(TokenType::IF);

    // Parse head
    this.parseAssignExpr();

    // Parse stmtLst
    this.parseStmtLst();

    // Parse else
    if !this.currentTokenIs(TokenType::ELSE) {
        this.parseElseStmt();
    }

    return this.concludeNode(ifStmtNode);
}

f<ASTElseStmtNode*> Parser.parseElseStmt() {
    dyn elseStmtNode = this.createNode<ASTElseStmtNode>();

    this.lexer.expect(TokenType::ELSE);

    if this.currentTokenIs(TokenType::IF) { // Else if
        this.parseIfStmt();
    } else { // Else
        this.parseStmtLst();
    }

    return this.concludeNode(elseStmtNode);
}

f<ASTSwitchStmtNode*> Parser.parseSwitchStmt() {
    dyn switchStmtNode = this.createNode<ASTSwitchStmtNode>();

    this.lexer.expect(TokenType::SWITCH);
    this.parseAssignExpr();
    this.lexer.expect(TokenType::LBRACE);
    while !this.currentTokenIs(TokenType::RBRACE) {
        this.parseCaseBranch();
    }
    if this.currentTokenIs(TokenType::DEFAULT) {
        this.parseDefaultBranch();
    }
    this.lexer.expect(TokenType::RBRACE);

    return this.concludeNode(switchStmtNode);
}

f<ASTCaseBranchNode*> Parser.parseCaseBranch() {
    dyn caseBranchNode = this.createNode<ASTCaseBranchNode>();

    this.lexer.expect(TokenType::CASE);
    this.parseCaseConstant();
    while this.currentTokenIs(TokenType::COMMA) {
        this.lexer.expect(TokenType::COMMA);
        this.parseCaseConstant();
    }
    this.lexer.expect(TokenType::COLON);
    this.parseStmtLst();

    return this.concludeNode(caseBranchNode);
}

f<ASTDefaultBranchNode*> Parser.parseDefaultBranch() {
    dyn defaultBranchNode = this.createNode<ASTDefaultBranchNode>();

    this.lexer.expect(TokenType::DEFAULT);
    this.lexer.expect(TokenType::COLON);
    this.parseStmtLst();

    return this.concludeNode(defaultBranchNode);
}

f<ASTAnonymousBlockStmtNode*> Parser.parseAnonymousBlockStmt() {
    dyn anonymousBlockStmtNode = this.createNode<ASTAnonymousBlockStmtNode>();

    this.parseStmtLst();

    return this.concludeNode(anonymousBlockStmtNode);
}

f<ASTStmtLstNode*> Parser.parseStmtLst() {
    dyn stmtLstNode = this.createNode<ASTStmtLstNode>();

    while !this.currentTokenIs(TokenType::RBRACE) {
        this.parseStmt();
    }

    return this.concludeNode(stmtLstNode);
}

f<ASTTypeLstNode*> Parser.parseTypeLst() {
    dyn typeLstNode = this.createNode<ASTTypeLstNode>();

    this.parseDataType();
    while this.currentTokenIs(TokenType::COMMA) {
        this.lexer.expect(TokenType::COMMA);
        this.parseDataType();
    }

    return this.concludeNode(typeLstNode);
}

f<ASTTypeAltsLstNode*> Parser.parseTypeAltsLst() {
    dyn typeAltsLstNode = this.createNode<ASTTypeAltsLstNode>();

    this.parseDataType();
    while this.currentTokenIs(TokenType::BITWISE_OR) {
        this.lexer.expect(TokenType::BITWISE_OR);
        this.parseDataType();
    }

    return this.concludeNode(typeAltsLstNode);
}

f<ASTParamLstNode*> Parser.parseParamLst() {
    dyn paramLstNode = this.createNode<ASTParamLstNode>();

    this.parseDeclStmt();
    while this.currentTokenIs(TokenType::COMMA) {
        this.lexer.expect(TokenType::COMMA);
        this.parseDeclStmt();
    }

    return this.concludeNode(paramLstNode);
}

f<ASTArgLstNode*> Parser.parseArgLst() {
    dyn argLstNode = this.createNode<ASTArgLstNode>();

    this.parseAssignExpr();
    while this.currentTokenIs(TokenType::COMMA) {
        this.lexer.expect(TokenType::COMMA);
        this.parseAssignExpr();
    }

    return this.concludeNode(argLstNode);
}

f<ASTEnumItemLstNode*> Parser.parseEnumItemLst() {
    dyn enumItemLstNode = this.createNode<ASTEnumItemLstNode>();

    this.parseEnumItem();
    while this.currentTokenIs(TokenType::COMMA) {
        this.lexer.expect(TokenType::COMMA);
        this.parseEnumItem();
    }

    return this.concludeNode(enumItemLstNode);
}

f<ASTEnumItemNode*> Parser.parseEnumItem() {
    dyn enumItemNode = this.createNode<ASTEnumItemNode>();

    this.lexer.expect(TokenType::TYPE_IDENTIFIER);
    if this.currentTokenIs(TokenType::ASSIGN) {
        this.lexer.expect(TokenType::ASSIGN);
        this.lexer.expect(TokenType::INT_LIT);
    }

    return this.concludeNode(enumItemNode);
}

f<ASTFieldNode*> Parser.parseField() {
    dyn fieldNode = this.createNode<ASTFieldNode>();

    this.parseDataType();
    this.lexer.expect(TokenType::IDENTIFIER);

    if this.currentTokenIs(TokenType::ASSIGN) {
        this.lexer.expect(TokenType::ASSIGN);
        this.parseTernaryExpr();
    }

    return this.concludeNode(fieldNode);
}

f<ASTSignatureNode*> Parser.parseSignature() {
    dyn signatureNode = this.createNode<ASTSignatureNode>();

    // Parse specifierLst
    const dyn options = [TokenType::F, TokenType::P];
    if !this.currentTokenIsOneOf(options, sizeof(options)) {
        this.parseSpecifierLst();
    }

    if this.currentTokenIs(TokenType::F) {
        this.lexer.expect(TokenType::F);
        this.lexer.expect(TokenType::LESS);
        this.parseDataType();
        this.lexer.expect(TokenType::GREATER);
    } else {
        this.lexer.expect(TokenType::P);
    }

    // Parse function name
    this.lexer.expect(TokenType::IDENTIFIER);

    // Parse typeLst (template type list)
    if this.currentTokenIs(TokenType::LESS) {
        this.lexer.expect(TokenType::LESS);
        this.parseTypeLst();
        this.lexer.expect(TokenType::GREATER);
    }

    // Parse paramLst
    this.lexer.expect(TokenType::LPAREN);
    if !this.currentTokenIs(TokenType::RPAREN) {
        this.parseParamLst();
    }
    this.lexer.expect(TokenType::RPAREN);

    this.lexer.expect(TokenType::SEMICOLON);

    return this.concludeNode(signatureNode);
}

f<ASTStmtNode*> Parser.parseStmt() {
    dyn stmtNode = this.createNode<ASTStmtNode>();

    const dyn declStmtSelect = [
        // declStmt -> dataType -> specifierLst -> specifier
        TokenType::CONST,
        TokenType::SIGNED,
        TokenType::UNSIGNED,
        TokenType::INLINE,
        TokenType::PUBLIC,
        TokenType::HEAP,
        TokenType::COMPOSE,
        // declStmt -> dataType -> baseDataType
        TokenType::TYPE_DOUBLE,
        TokenType::TYPE_INT,
        TokenType::TYPE_SHORT,
        TokenType::TYPE_LONG,
        TokenType::TYPE_BYTE,
        TokenType::TYPE_CHAR,
        TokenType::TYPE_STRING,
        TokenType::TYPE_BOOL,
        TokenType::TYPE_DYN
        // ToDo: add other
    ];
    if this.currentTokenIs(TokenType::RETURN) {
        this.parseReturnStmt();
    } else if this.currentTokenIs(TokenType::BREAK) {
        this.parseBreakStmt();
    } else if this.currentTokenIs(TokenType::CONTINUE) {
        this.parseContinueStmt();
    } else if this.currentTokenIs(TokenType::FALLTHROUGH) {
        this.parseFallthroughStmt();
    } else if this.currentTokenIsOneOf(declStmtSelect, sizeof(declStmtSelect)) {
        this.parseDeclStmt();
    } else {
        this.parseAssignExpr();
    }
    this.lexer.expect(TokenType::SEMICOLON);

    return this.concludeNode(stmtNode);
}

f<ASTDeclStmtNode*> Parser.parseDeclStmt() {
    dyn declStmtNode = this.createNode<ASTDeclStmtNode>();

    // Parse dataType
    this.parseDataType();

    this.lexer.expect(TokenType::IDENTIFIER);

    // Parse initializer
    if this.currentTokenIs(TokenType::ASSIGN) {
        this.lexer.expect(TokenType::ASSIGN);
        this.parseAssignExpr();
    }

    return this.concludeNode(declStmtNode);
}

f<ASTSpecifierLstNode*> Parser.parseSpecifierLst() {
    dyn specifierLstNode = this.createNode<ASTSpecifierLstNode>();

    const dyn specifierSelect = [TokenType::CONST, TokenType::SIGNED, TokenType::UNSIGNED, TokenType::INLINE, TokenType::PUBLIC, TokenType::HEAP, TokenType::COMPOSE];
    do {
        this.parseSpecifier();
    } while this.currentTokenIsOneOf(specifierSelect, sizeof(specifierSelect));

    return this.concludeNode(specifierLstNode);
}

f<ASTSpecifierNode*> Parser.parseSpecifier() {
    dyn specifierNode = this.createNode<ASTSpecifierNode>();

    if this.currentTokenIs(TokenType::CONST) {
        specifierNode.specifierType = SpecifierType::CONST;
    } else if this.currentTokenIs(TokenType::SIGNED) {
        specifierNode.specifierType = SpecifierType::SIGNED;
    } else if this.currentTokenIs(TokenType::UNSIGNED) {
        specifierNode.specifierType = SpecifierType::UNSIGNED;
    } else if this.currentTokenIs(TokenType::INLINE) {
        specifierNode.specifierType = SpecifierType::INLINE;
    } else if this.currentTokenIs(TokenType::PUBLIC) {
        specifierNode.specifierType = SpecifierType::PUBLIC;
    } else if this.currentTokenIs(TokenType::HEAP) {
        specifierNode.specifierType = SpecifierType::HEAP;
    } else if this.currentTokenIs(TokenType::COMPOSE) {
        specifierNode.specifierType = SpecifierType::COMPOSE;
    } else {
        assert false;
    }

    return this.concludeNode(specifierNode);
}

f<ASTModAttrNode*> Parser.parseModAttr() {
    dyn modAttrNode = this.createNode<ASTModAttrNode>();

    this.lexer.expect(TokenType::MOD_ATTR_PREAMBLE);
    this.lexer.expect(TokenType::LBRACKET);
    this.parseAttrLst();
    this.lexer.expect(TokenType::RBRACKET);

    return this.concludeNode(modAttrNode);
}

f<ASTTopLevelDefAttrNode*> Parser.parseTopLevelDefAttr() {
    dyn topLevelDefAttrNode = this.createNode<ASTTopLevelDefAttrNode>();

    this.lexer.expect(TokenType::FCT_ATTR_PREAMBLE);
    this.lexer.expect(TokenType::LBRACKET);
    this.parseAttrLst();
    this.lexer.expect(TokenType::RBRACKET);

    return this.concludeNode(topLevelDefAttrNode);
}

f<ASTLambdaAttrNode*> Parser.parseLambdaAttr() {
    dyn lambdaAttrNode = this.createNode<ASTLambdaAttrNode>();

    this.lexer.expect(TokenType::LBRACKET);
    this.lexer.expect(TokenType::LBRACKET);
    this.parseAttrLst();
    this.lexer.expect(TokenType::RBRACKET);
    this.lexer.expect(TokenType::RBRACKET);

    return this.concludeNode(lambdaAttrNode);
}

f<ASTAttrLstNode*> Parser.parseAttrLst() {
    dyn attrLstNode = this.createNode<ASTAttrLstNode>();

    this.parseAttr();
    while this.currentTokenIs(TokenType::COMMA) {
        this.lexer.expect(TokenType::COMMA);
        this.parseAttr();
    }

    return this.concludeNode(attrLstNode);
}

f<ASTAttrNode*> Parser.parseAttr() {
    dyn attrNode = this.createNode<ASTAttrNode>();

    // Parse attribute name
    this.lexer.expect(TokenType::IDENTIFIER);
    while this.currentTokenIs(TokenType::DOT) {
        this.lexer.expect(TokenType::DOT);
        this.lexer.expect(TokenType::IDENTIFIER);
    }

    // Parse attribute value
    if this.currentTokenIs(TokenType::ASSIGN) {
        this.lexer.expect(TokenType::ASSIGN);
        this.parseConstant();
    }

    return this.concludeNode(attrNode);
}

f<ASTCaseConstantNode*> Parser.parseCaseConstant() {
    dyn caseConstantNode = this.createNode<ASTCaseConstantNode>();

    const dyn optionsVarExpr = [TokenType::IDENTIFIER, TokenType::TYPE_IDENTIFIER];
    if this.currentTokenIsOneOf(optionsVarExpr, sizeof(optionsVarExpr)) {
        if this.currentTokenIs(TokenType::TYPE_IDENTIFIER) {
            this.lexer.advance();
            this.lexer.expect(TokenType::SCOPE_ACCESS);
        }
        this.lexer.expect(TokenType::TYPE_IDENTIFIER);
        while this.currentTokenIs(TokenType::SCOPE_ACCESS) {
            this.lexer.expect(TokenType::SCOPE_ACCESS);
            this.lexer.expect(TokenType::TYPE_IDENTIFIER);
        }
    } else {
        this.parseConstant();
    }

    return this.concludeNode(caseConstantNode);
}

f<ASTReturnStmtNode*> Parser.parseReturnStmt() {
    dyn returnStmtNode = this.createNode<ASTReturnStmtNode>();

    this.lexer.expect(TokenType::RETURN);
    if !this.currentTokenIs(TokenType::SEMICOLON) {
        this.parseAssignExpr();
    }

    return this.concludeNode(returnStmtNode);
}

f<ASTBreakStmtNode*> Parser.parseBreakStmt() {
    dyn breakStmtNode = this.createNode<ASTBreakStmtNode>();

    this.lexer.expect(TokenType::BREAK);
    if this.currentTokenIs(TokenType::INT_LIT) {
        this.lexer.expect(TokenType::INT_LIT);
    }

    return this.concludeNode(breakStmtNode);
}

f<ASTContinueStmtNode*> Parser.parseContinueStmt() {
    dyn continueStmtNode = this.createNode<ASTContinueStmtNode>();

    this.lexer.expect(TokenType::CONTINUE);
    if this.currentTokenIs(TokenType::INT_LIT) {
        this.lexer.expect(TokenType::INT_LIT);
    }

    return this.concludeNode(continueStmtNode);
}

f<ASTFallthroughStmtNode*> Parser.parseFallthroughStmt() {
    dyn fallthroughStmtNode = this.createNode<ASTFallthroughStmtNode>();

    this.lexer.expect(TokenType::FALLTHROUGH);

    return this.concludeNode(fallthroughStmtNode);
}

f<ASTAssertStmtNode*> Parser.parseAssertStmt() {
    dyn assertStmtNode = this.createNode<ASTAssertStmtNode>();

    this.lexer.expect(TokenType::ASSERT);
    this.parseAssignExpr();
    this.lexer.expect(TokenType::SEMICOLON);

    return this.concludeNode(assertStmtNode);
}

f<ASTPrintfCallNode*> Parser.parsePrintfCall() {
    dyn printfCallNode = this.createNode<ASTPrintfCallNode>();

    this.lexer.expect(TokenType::PRINTF);
    this.lexer.expect(TokenType::LPAREN);
    this.lexer.expect(TokenType::STRING_LIT);
    while this.currentTokenIs(TokenType::COMMA) {
        this.lexer.expect(TokenType::COMMA);
        this.parseAssignExpr();
    }
    this.lexer.expect(TokenType::RPAREN);

    return this.concludeNode(printfCallNode);
}

f<ASTSizeofCallNode*> Parser.parseSizeOfCall() {
    dyn sizeofCallNode = this.createNode<ASTSizeofCallNode>();

    this.lexer.expect(TokenType::SIZEOF);
    this.lexer.expect(TokenType::LPAREN);

    if this.currentTokenIs(TokenType::TYPE) {
        this.lexer.expect(TokenType::TYPE);
        this.parseDataType();
    } else {
        this.parseAssignExpr();
    }

    this.lexer.expect(TokenType::RPAREN);

    return this.concludeNode(sizeofCallNode);
}

f<ASTAlignofCallNode*> Parser.parseAlignOfCall() {
    dyn alignofCallNode = this.createNode<ASTAlignofCallNode>();

    this.lexer.expect(TokenType::ALIGNOF);
    this.lexer.expect(TokenType::LPAREN);

    if this.currentTokenIs(TokenType::TYPE) {
        this.lexer.expect(TokenType::TYPE);
        this.parseDataType();
    } else {
        this.parseAssignExpr();
    }

    this.lexer.expect(TokenType::RPAREN);

    return this.concludeNode(alignofCallNode);
}

f<ASTLenCallNode*> Parser.parseLenCall() {
    dyn lenCallNode = this.createNode<ASTLenCallNode>();

    this.lexer.expect(TokenType::LEN);
    this.lexer.expect(TokenType::LPAREN);
    this.parseAssignExpr();
    this.lexer.expect(TokenType::RPAREN);

    return this.concludeNode(lenCallNode);
}

f<ASTPanicCallNode*> Parser.parsePanicCall() {
    dyn panicCallNode = this.createNode<ASTPanicCallNode>();

    this.lexer.expect(TokenType::PANIC);
    this.lexer.expect(TokenType::LPAREN);
    this.parseAssignExpr();
    this.lexer.expect(TokenType::RPAREN);

    return this.concludeNode(panicCallNode);
}

f<ASTAssignExprNode*> Parser.parseAssignExpr() {
    dyn assignExprNode = this.createNode<ASTAssignExprNode>();

    // ToDo: implement

    return this.concludeNode(assignExprNode);
}

f<ASTTernaryExprNode*> Parser.parseTernaryExpr() {
    dyn ternaryExprNode = this.createNode<ASTTernaryExprNode>();

    // Parse lhs
    this.parseLogicalOrExpr();

    // Parse both rhs branches
    if this.currentTokenIs(TokenType::QUESTION_MARK) {
        this.lexer.expect(TokenType::QUESTION_MARK);
        this.parseLogicalOrExpr();
        this.lexer.expect(TokenType::COLON);
        this.parseLogicalOrExpr();
    }

    return this.concludeNode(ternaryExprNode);
}

f<ASTLogicalOrExprNode*> Parser.parseLogicalOrExpr() {
    dyn logicalOrExprNode = this.createNode<ASTLogicalOrExprNode>();

    // Parse lhs
    this.parseLogicalAndExpr();

    // Parse rhs
    while this.currentTokenIs(TokenType::LOGICAL_OR) {
        this.lexer.expect(TokenType::LOGICAL_OR);
        this.parseLogicalAndExpr();
    }

    return this.concludeNode(logicalOrExprNode);
}

f<ASTLogicalAndExprNode*> Parser.parseLogicalAndExpr() {
    dyn logicalAndExprNode = this.createNode<ASTLogicalAndExprNode>();

    // Parse lhs
    this.parseBitwiseOrExpr();

    // Parse rhs
    while this.currentTokenIs(TokenType::LOGICAL_AND) {
        this.lexer.expect(TokenType::LOGICAL_AND);
        this.parseBitwiseOrExpr();
    }

    return this.concludeNode(logicalAndExprNode);
}

f<ASTBitwiseOrExprNode*> Parser.parseBitwiseOrExpr() {
    dyn bitwiseOrExprNode = this.createNode<ASTBitwiseOrExprNode>();

    // Parse lhs
    this.parseBitwiseXorExpr();

    // Parse rhs
    while this.currentTokenIs(TokenType::BITWISE_OR) {
        this.lexer.expect(TokenType::BITWISE_OR);
        this.parseBitwiseXorExpr();
    }

    return this.concludeNode(bitwiseOrExprNode);
}

f<ASTBitwiseXorExprNode*> Parser.parseBitwiseXorExpr() {
    dyn bitwiseXorExprNode = this.createNode<ASTBitwiseXorExprNode>();

    // Parse lhs
    this.parseBitwiseAndExpr();

    // Parse rhs
    while this.currentTokenIs(TokenType::BITWISE_XOR) {
        this.lexer.expect(TokenType::BITWISE_XOR);
        this.parseBitwiseAndExpr();
    }

    return this.concludeNode(bitwiseXorExprNode);
}

f<ASTBitwiseAndExprNode*> Parser.parseBitwiseAndExpr() {
    dyn bitwiseAndExprNode = this.createNode<ASTBitwiseAndExprNode>();

    // Parse lhs
    this.parseEqualityExpr();

    // Parse rhs
    while this.currentTokenIs(TokenType::BITWISE_AND) {
        this.lexer.expect(TokenType::BITWISE_AND);
        this.parseEqualityExpr();
    }

    return this.concludeNode(bitwiseAndExprNode);
}

f<ASTEqualityExprNode*> Parser.parseEqualityExpr() {
    dyn equalityExprNode = this.createNode<ASTEqualityExprNode>();

    // Parse lhs
    this.parseRelationalExpr();

    // Parse rhs
    const dyn options = [TokenType::EQUAL, TokenType::NOT_EQUAL];
    while this.currentTokenIsOneOf(options, sizeof(options)) {
        this.lexer.advance();
        this.parseRelationalExpr();
    }

    return this.concludeNode(equalityExprNode);
}

f<ASTRelationalExprNode*> Parser.parseRelationalExpr() {
    dyn relationalExprNode = this.createNode<ASTRelationalExprNode>();

    // Parse lhs
    this.parseShiftExpr();

    // Parse rhs
    const dyn optionsRelationalOp = [TokenType::LESS, TokenType::GREATER, TokenType::LESS_EQUAL, TokenType::GREATER_EQUAL];
    while this.currentTokenIsOneOf(optionsRelationalOp, sizeof(optionsRelationalOp)) {
        this.lexer.advance();
        this.parseShiftExpr();
    }

    return this.concludeNode(relationalExprNode);
}

f<ASTShiftExprNode*> Parser.parseShiftExpr() {
    dyn shiftExprNode = this.createNode<ASTShiftExprNode>();

    // Parse lhs
    this.parseAdditiveExpr();

    // Parse rhs
    const dyn options = [TokenType::LESS, TokenType::GREATER];
    while this.currentTokenIsOneOf(options, sizeof(options)) {
        this.lexer.advance();
        assert this.currentTokenIsOneOf(options, sizeof(options));
        this.lexer.advance();
        this.parseAdditiveExpr();
    }

    return this.concludeNode(shiftExprNode);
}

f<ASTAdditiveExprNode*> Parser.parseAdditiveExpr() {
    dyn additiveExprNode = this.createNode<ASTAdditiveExprNode>();

    // Parse lhs
    this.parseMultiplicativeExpr();

    // Parse rhs
    const dyn options = [TokenType::PLUS, TokenType::MINUS];
    while this.currentTokenIsOneOf(options, sizeof(options)) {
        this.lexer.advance();
        this.parseMultiplicativeExpr();
    }

    return this.concludeNode(additiveExprNode);
}

f<ASTMultiplicativeExprNode*> Parser.parseMultiplicativeExpr() {
    dyn multiplicativeExprNode = this.createNode<ASTMultiplicativeExprNode>();

    // Parse lhs
    this.parseCastExpr();

    // Parse rhs
    const dyn options = [TokenType::MUL, TokenType::DIV, TokenType::REM];
    while this.currentTokenIsOneOf(options, sizeof(options)) {
        this.lexer.advance();
        this.parseCastExpr();
    }

    return this.concludeNode(multiplicativeExprNode);
}

f<ASTCastExprNode*> Parser.parseCastExpr() {
    dyn castExprNode = this.createNode<ASTCastExprNode>();

    // Parse target type
    this.lexer.expect(TokenType::LPAREN);
    this.parseDataType();
    this.lexer.expect(TokenType::RPAREN);

    // Parse rhs
    this.parsePrefixUnaryExpr();

    return this.concludeNode(castExprNode);
}

f<ASTPrefixUnaryExprNode*> Parser.parsePrefixUnaryExpr() {
    dyn prefixUnaryExprNode = this.createNode<ASTPrefixUnaryExprNode>();

    const dyn options = [TokenType::MINUS, TokenType::PLUS_PLUS, TokenType::MINUS_MINUS, TokenType::NOT, TokenType::BITWISE_NOT, TokenType::MUL, TokenType::BITWISE_AND];
    if this.currentTokenIsOneOf(options, sizeof(options)) {
        this.lexer.advance();
        this.parsePrefixUnaryExpr();
    } else {
        this.parsePostfixUnaryExpr();
    }

    return this.concludeNode(prefixUnaryExprNode);
}

f<ASTPostfixUnaryExprNode*> Parser.parsePostfixUnaryExpr() {
    dyn postfixUnaryExprNode = this.createNode<ASTPostfixUnaryExprNode>();

    // ToDo: Implement

    return this.concludeNode(postfixUnaryExprNode);
}

f<ASTAtomicExprNode*> Parser.parseAtomicExpr() {
    dyn atomicExprNode = this.createNode<ASTAtomicExprNode>();

    const dyn optionsVarExpr = [TokenType::IDENTIFIER, TokenType::TYPE_IDENTIFIER];
    const dyn optionsConstant = [TokenType::DOUBLE_LIT, TokenType::INT_LIT, TokenType::SHORT_LIT, TokenType::LONG_LIT, TokenType::CHAR_LIT, TokenType::STRING_LIT, TokenType::TRUE, TokenType::FALSE];

    if this.currentTokenIsOneOf(optionsVarExpr, sizeof(optionsVarExpr)) {
        this.lexer.advance();
        while this.currentTokenIs(TokenType::SCOPE_ACCESS) {
            this.lexer.expect(TokenType::SCOPE_ACCESS);
            if this.currentTokenIs(TokenType::TYPE_IDENTIFIER) {
                this.lexer.expect(TokenType::TYPE_IDENTIFIER);
            } else {
                this.lexer.expect(TokenType::IDENTIFIER);
            }
        }
    } else if this.currentTokenIsOneOf(optionsConstant, sizeof(optionsConstant)) {
        this.parseConstant();
    } else if this.currentTokenIs(TokenType::PRINTF) {
        this.parsePrintfCall();
    } else if this.currentTokenIs(TokenType::SIZEOF) {
        this.parseSizeOfCall();
    } else if this.currentTokenIs(TokenType::ALIGNOF) {
        this.parseAlignOfCall();
    } else if this.currentTokenIs(TokenType::LEN) {
        this.parseLenCall();
    } else if this.currentTokenIs(TokenType::PANIC) {
        this.parsePanicCall();
    } else if this.currentTokenIs(TokenType::LPAREN) {
        this.lexer.expect(TokenType::LPAREN);
        this.parseAssignExpr();
        this.lexer.expect(TokenType::RPAREN);
    } else {
        this.parseValue();
    }

    return this.concludeNode(atomicExprNode);
}

f<ASTValueNode*> Parser.parseValue() {
    dyn valueNode = this.createNode<ASTValueNode>();

    // ToDo: Implement

    return this.concludeNode(valueNode);
}

f<ASTConstantNode*> Parser.parseConstant() {
    dyn constantNode = this.createNode<ASTConstantNode>();

    // ToDo: Implement

    return this.concludeNode(constantNode);
}

f<ASTFctCallNode*> Parser.parseFctCall() {
    dyn fctCallNode = this.createNode<ASTFctCallNode>();

    // ToDo: Implement

    return this.concludeNode(fctCallNode);
}

f<ASTArrayInitializationNode*> Parser.parseArrayInitialization() {
    dyn arrayInitializationNode = this.createNode<ASTArrayInitializationNode>();

    this.lexer.expect(TokenType::LBRACKET);
    this.parseArgLst();
    this.lexer.expect(TokenType::RBRACKET);

    return this.concludeNode(arrayInitializationNode);
}

f<ASTStructInstantiationNode*> Parser.parseStructInstantiation() {
    dyn structInstantiationNode = this.createNode<ASTStructInstantiationNode>();

    while !this.currentTokenIs(TokenType::IDENTIFIER) {
        this.lexer.expect(TokenType::IDENTIFIER);
        this.lexer.expect(TokenType::SCOPE_ACCESS);
    }

    this.lexer.expect(TokenType::TYPE_IDENTIFIER);

    if this.currentTokenIs(TokenType::LESS) {
        this.lexer.expect(TokenType::LESS);
        this.parseTypeLst();
        this.lexer.expect(TokenType::GREATER);
    }

    this.lexer.expect(TokenType::LBRACE);
    this.parseArgLst();
    this.lexer.expect(TokenType::RBRACE);

    return this.concludeNode(structInstantiationNode);
}

f<ASTLambdaFuncNode*> Parser.parseLambdaFunc() {
    dyn lambdaFuncNode = this.createNode<ASTLambdaFuncNode>();

    this.lexer.expect(TokenType::F);
    this.lexer.expect(TokenType::LESS);
    this.parseDataType();
    this.lexer.expect(TokenType::GREATER);
    this.lexer.expect(TokenType::LPAREN);
    if !this.currentTokenIs(TokenType::RPAREN) {
        this.parseParamLst();
    }
    this.lexer.expect(TokenType::RPAREN);

    // Parse lambda attrs
    if this.currentTokenIs(TokenType::LBRACKET) {
        this.parseLambdaAttr();
    }

    this.parseStmtLst();

    return this.concludeNode(lambdaFuncNode);
}

f<ASTLambdaProcNode*> Parser.parseLambdaProc() {
    dyn lambdaProcNode = this.createNode<ASTLambdaProcNode>();

    this.lexer.expect(TokenType::P);

    // Parse paramLst
    this.lexer.expect(TokenType::LPAREN);
    if !this.currentTokenIs(TokenType::RPAREN) {
        this.parseParamLst();
    }
    this.lexer.expect(TokenType::RPAREN);

    // Parse lambda attrs
    if this.currentTokenIs(TokenType::LBRACKET) {
        this.parseLambdaAttr();
    }

    // Parse
    this.parseStmtLst();

    return this.concludeNode(lambdaProcNode);
}

f<ASTLambdaExprNode*> Parser.parseLambdaExpr() {
    dyn lambdaExprNode = this.createNode<ASTLambdaExprNode>();

    // Parse paramLst
    this.lexer.expect(TokenType::LPAREN);
    if !this.currentTokenIs(TokenType::RPAREN) {
        this.parseParamLst();
    }
    this.lexer.expect(TokenType::RPAREN);

    this.lexer.expect(TokenType::ARROW);
    this.parseAssignExpr();

    return this.concludeNode(lambdaExprNode);
}

f<ASTDataTypeNode*> Parser.parseDataType() {
    dyn dataTypeNode = this.createNode<ASTDataTypeNode>();

    const dyn optionsSpecifierLst = [TokenType::CONST, TokenType::SIGNED, TokenType::UNSIGNED, TokenType::INLINE, TokenType::PUBLIC, TokenType::HEAP, TokenType::COMPOSE];
    if this.currentTokenIsOneOf(optionsSpecifierLst, sizeof(optionsSpecifierLst)) {
        this.parseSpecifierLst();
    }
    this.parseBaseDataType();

    // ToDo: Implement

    return this.concludeNode(dataTypeNode);
}

f<ASTBaseDataTypeNode*> Parser.parseBaseDataType() {
    dyn baseDataTypeNode = this.createNode<ASTBaseDataTypeNode>();

    const dyn optionsFctDataType = [TokenType::F, TokenType::P];
    if this.currentTokenIs(TokenType::TYPE_DOUBLE) {
        this.lexer.expect(TokenType::TYPE_DOUBLE);
    } else if this.currentTokenIs(TokenType::TYPE_INT) {
        this.lexer.expect(TokenType::TYPE_INT);
    } else if this.currentTokenIs(TokenType::TYPE_SHORT) {
        this.lexer.expect(TokenType::TYPE_SHORT);
    } else if this.currentTokenIs(TokenType::TYPE_LONG) {
        this.lexer.expect(TokenType::TYPE_LONG);
    } else if this.currentTokenIs(TokenType::TYPE_BYTE) {
        this.lexer.expect(TokenType::TYPE_BYTE);
    } else if this.currentTokenIs(TokenType::TYPE_CHAR) {
        this.lexer.expect(TokenType::TYPE_CHAR);
    } else if this.currentTokenIs(TokenType::TYPE_STRING) {
        this.lexer.expect(TokenType::TYPE_STRING);
    } else if this.currentTokenIs(TokenType::TYPE_BOOL) {
        this.lexer.expect(TokenType::TYPE_BOOL);
    } else if this.currentTokenIs(TokenType::TYPE_DYN) {
        this.lexer.expect(TokenType::TYPE_DYN);
    } else if this.currentTokenIsOneOf(optionsFctDataType, sizeof(optionsFctDataType)) {
        this.parseFunctionDataType();
    } else {
        this.parseCustomDataType();
    }

    return this.concludeNode(baseDataTypeNode);
}

f<ASTCustomDataTypeNode*> Parser.parseCustomDataType() {
    dyn customDataTypeNode = this.createNode<ASTCustomDataTypeNode>();

    // Parse type name
    while !this.currentTokenIs(TokenType::TYPE_IDENTIFIER) {
        this.lexer.expect(TokenType::IDENTIFIER);
        this.lexer.expect(TokenType::SCOPE_ACCESS);
    }
    this.lexer.expect(TokenType::TYPE_IDENTIFIER);

    // Parse typeLst (template type list)
    if this.currentTokenIs(TokenType::LESS) {
        this.lexer.expect(TokenType::LESS);
        this.parseTypeLst();
        this.lexer.expect(TokenType::GREATER);
    }

    return this.concludeNode(customDataTypeNode);
}

f<ASTFunctionDataTypeNode*> Parser.parseFunctionDataType() {
    dyn functionDataTypeNode = this.createNode<ASTFunctionDataTypeNode>();

    if this.currentTokenIs(TokenType::F) {
        this.lexer.expect(TokenType::F);
        this.lexer.expect(TokenType::LESS);
        this.parseDataType();
        this.lexer.expect(TokenType::GREATER);
    } else {
        this.lexer.expect(TokenType::P);
    }

    // Parse typeLst (param types)
    this.lexer.expect(TokenType::LPAREN);
    if !this.currentTokenIs(TokenType::RPAREN) {
        this.parseTypeLst();
    }
    this.lexer.expect(TokenType::RPAREN);

    return this.concludeNode(functionDataTypeNode);
}