// Std imports
import "std/io/filepath";
import "std/io/file";
import "std/type/result";
import "std/type/error";
import "std/os/os";

// Own imports
import "../reader/code-loc";

public type Reader struct {
    File file
    string filename
    char curChar = '\0'
    CodeLoc curCodeLoc
}

public p Reader.ctor(string inputFileName) {
    this.filename = inputFileName;
    this.curCodeLoc = CodeLoc(1l, 0l, inputFileName);

    // Open the file input stream
    Result<File> result = openFile(inputFileName, MODE_READ);
    if !result.isOk() {
        panic(Error("Source file cannot be opened"));
    }
    this.file = result.unwrap();

    // Read the first character
    this.advance();
}

/**
 * Get the previously read character
 *
 * @return char Last character
 */
public inline f<char> Reader.getChar() {
    return this.curChar;
}

/**
 * Get the code location of the previously read character
 *
 * @return CodeLoc Code location
 */
public inline f<CodeLoc&> Reader.getCodeLoc() {
    return this.curCodeLoc;
}

/**
 * Advance the reader by one character
 */
public p Reader.advance() {
    assert !this.isEOF();
    this.curChar = this.file.readChar();
    if this.curChar == '\n' {
        this.curCodeLoc.line++;
        this.curCodeLoc.col = 0l;
    }
    this.curCodeLoc.col++;
}

/**
 * Advance the reader by one character and check if this char equals the expected.
 *
 * @param c Expected char
 */
public inline p Reader.expect(char c) {
    assert this.curChar == c;
    this.advance();
}

/**
 * Check if we are at the end of the input file
 *
 * @return At the end or not
 */
public inline f<bool> Reader.isEOF() {
    return this.file.isEOF();
}