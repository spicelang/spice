public const int SIZE = 32;
public const int MIN_VALUE = -2147483648;
public const int MAX_VALUE = 2147483647;

// Converts an int to a double
public f<double> toDouble(int input) {
    // ToDo: Implement
    return 0.0;
}

// Converts an int to a short
public f<short> toShort(int input) {
    return (short) input;
}

// Converts an int to a long
public f<long> toLong(int input) {
    return (long) input;
}

// Converts an int to a byte
public f<byte> toByte(int input) {
    return (byte) input;
}

// Converts an int to a char
public f<char> toChar(int input) {
    return (char) input;
}

// Converts an int to a string
public f<string> toString(int input) {
    // ToDo: Implement (See https://github.com/golang/go/blob/master/src/strconv/itoa.go)
    return "";
}

// Converts an int to a boolean
public f<bool> toBool(int input) {
    return input >= 1;
}