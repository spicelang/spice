f<bool> fn(int& ref) {
    return false;
}

f<int> main() {
    fn(123);
}