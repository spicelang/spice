import "std/data/optional";
import "std/data/stack";

f<int> main() {
    Stack<double> doubleStack = Stack<double>();
    doubleStack.push(4.566);

    dyn oi = Optional<Stack<double>>();
    printf("%d\n", oi.isPresent());
    oi.set(doubleStack);
    printf("%d\n", oi.isPresent());
    printf("%d\n", oi.get().getSize());
    oi.clear();
    printf("%d\n", oi.isPresent());
    assert oi.get() == nil<Stack<double>>;
}