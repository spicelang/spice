f<int> main() {
    int t = 123;
    heap int* test = &t;
}