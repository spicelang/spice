f<int> main() {
    
}