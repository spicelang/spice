f<int> getAge() {
    dyn i;
    bool b = true;
    if (b) {
        result = 20;
        return;
    } else if (i = false) {
        result = 19;
    }
    result = 18;
}

f<int> main() {
    int age = getAge();
    printf("The age is: %d", age);
}