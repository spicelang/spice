f<int> main() {
    int variable = 12;
    if (true) {
        variable++;
        double variable = 14.1;
        printf("Inner variable: %f\n", variable);
    }
    printf("Outer variable: %d", variable);
}