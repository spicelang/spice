// Converts an integer to a double
f<double> toDouble(int number) {
    return number + 0.0;
}

// Converts a string to a double
f<double> toDouble(string text) {
    return 0.0; // ToDo: not implemented
}

// Converts a double to an integer
f<int> toInt(double fp) {
    return 0; // ToDo: not implemented
}

// Converts a string to an integer
f<int> toInt(string text) {
    return 0; // ToDo: not implemented
}

// Converts a boolean to an integer
f<int> toInt(bool value) {
    return value ? 1 : 0;
}

// Converts a double to a string
f<string> toString(double number) {
    return "0.0"; // ToDo: not implemented
}

// Converts an integer to a string
f<string> toString(int number) {
    return "0"; // ToDo: not implemented
}

// Converts a boolean to a string
f<string> toString(bool value) {
    return value ? "true" : "false";
}

/*// Converts a double to a bool
f<bool> toString(double number) {
    return number >= 0.5 ? true : false;
}

// Converts an integer to a bool
f<bool> toString(int number) {
    return number > 0 ? true : false;
}

// Converts a string to a bool
f<bool> toString(string text) {
    return text == "true" ? true : false;
}*/