f<int> main() {
    int test = 123;
    int& testRef = test;
    assert &test == &testRef;
}