import "std/runtime/iterator_rt";

f<int> main() {
    // Create test array to iterate over
    int[5] a = { 123, 4321, 9876, 321, -99 };

    foreach int& aItem : iterate(a, len(a)) {
        printf("%d\n", aItem);
    }

    printf("All assertions passed!");
}