// Common type aliases
type Size alias long;