import "std/test/assertions";

f<int> main() {
    assertTrue(2 != 1);
    assertFalse(7 == 1);
    assertEqual(6, 1 + 5);
    assertEqual("expected", false ? "actual" : "expected");
    assertNotEqual(7, 5 + 1);
    assertNil(nil<int>);
    assertNotNil(764s);
    assertEmpty("");
    assertNotEmpty("This is not an empty string");
    assertContains("This haystack contains some needles.", "needle");
    printf("All assertions passed!");
}