import "std/type/bool" as boolTy;

f<int> main() {
    printf("Result: %d\n", toInt(true));
}