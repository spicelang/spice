f<int> main() {
    f<int>(bool&) si = f<int>(bool& input) {
        if (!input) {
            input = false;
        } else {
            return 2;
        }
    };
    si(false);
}