#![
    // Paths - Linux
    core.linux.linker.flag = "-L$LLVM_LIB_DIR",
    core.linux.linker.flag = "-I$LLVM_INCLUDE_DIR",
    core.linux.linker.flag = "-I$LLVM_BUILD_INCLUDE_DIR",
    core.linux.linker.flag = "-lm", // math
    core.linux.linker.flag = "-lz", // zlib
    core.linux.linker.flag = "-ltinfo", // ncurses
    core.linux.linker.flag = "-lzstd", // zstd
    core.linux.linker.flag = "-luuid", // uuid
    // Paths - macOS
    core.darwin.linker.flag = "-L$LLVM_LIB_DIR",
    core.darwin.linker.flag = "-I$LLVM_INCLUDE_DIR",
    core.darwin.linker.flag = "-I$LLVM_BUILD_INCLUDE_DIR",
    core.darwin.linker.flag = "-lm", // math
    core.darwin.linker.flag = "-lz", // zlib
    core.darwin.linker.flag = "-lncurses", // ncurses
    core.darwin.linker.flag = "-lzstd", // zstd
    // Paths - Windows
    core.windows.linker.flag = "-L%LLVM_LIB_DIR%",           // e.g.: D:/LLVM/build-release/lib
    core.windows.linker.flag = "-I%LLVM_INCLUDE_DIR%",       // e.g.: D:/LLVM/llvm/include
    core.windows.linker.flag = "-I%LLVM_BUILD_INCLUDE_DIR%", // e.g.: D:/LLVM/build-release/include
    // Additional libs for Windows (taken from llvm/lib/Support/CMakeLists.txt)
    core.windows.linker.flag = "-lole32", // COM
    core.windows.linker.flag = "-lws2_32", // WinSock
    core.windows.linker.flag = "-lntdll", // Low level functions like syscalls
    core.windows.linker.flag = "-luuid", // uuid
    // LLVM libs
    core.linker.flag = "-lLLVMAArch64AsmParser",
    core.linker.flag = "-lLLVMAArch64CodeGen",
    core.linker.flag = "-lLLVMAArch64Desc",
    core.linker.flag = "-lLLVMAArch64Disassembler",
    core.linker.flag = "-lLLVMAArch64Info",
    core.linker.flag = "-lLLVMAArch64Utils",
    core.linker.flag = "-lLLVMAggressiveInstCombine",
    core.linker.flag = "-lLLVMAMDGPUAsmParser",
    core.linker.flag = "-lLLVMAMDGPUCodeGen",
    core.linker.flag = "-lLLVMAMDGPUDesc",
    core.linker.flag = "-lLLVMAMDGPUDisassembler",
    core.linker.flag = "-lLLVMAMDGPUInfo",
    core.linker.flag = "-lLLVMAMDGPUTargetMCA",
    core.linker.flag = "-lLLVMAMDGPUUtils",
    core.linker.flag = "-lLLVMAnalysis",
    core.linker.flag = "-lLLVMARMAsmParser",
    core.linker.flag = "-lLLVMARMCodeGen",
    core.linker.flag = "-lLLVMARMDesc",
    core.linker.flag = "-lLLVMARMDisassembler",
    core.linker.flag = "-lLLVMARMInfo",
    core.linker.flag = "-lLLVMARMUtils",
    core.linker.flag = "-lLLVMAsmParser",
    core.linker.flag = "-lLLVMAsmPrinter",
    core.linker.flag = "-lLLVMAVRAsmParser",
    core.linker.flag = "-lLLVMAVRCodeGen",
    core.linker.flag = "-lLLVMAVRDesc",
    core.linker.flag = "-lLLVMAVRDisassembler",
    core.linker.flag = "-lLLVMAVRInfo",
    core.linker.flag = "-lLLVMBinaryFormat",
    core.linker.flag = "-lLLVMBitReader",
    core.linker.flag = "-lLLVMBitstreamReader",
    core.linker.flag = "-lLLVMBitWriter",
    core.linker.flag = "-lLLVMBPFAsmParser",
    core.linker.flag = "-lLLVMBPFCodeGen",
    core.linker.flag = "-lLLVMBPFDesc",
    core.linker.flag = "-lLLVMBPFDisassembler",
    core.linker.flag = "-lLLVMBPFInfo",
    core.linker.flag = "-lLLVMCFGuard",
    core.linker.flag = "-lLLVMCFIVerify",
    core.linker.flag = "-lLLVMCGData",
    core.linker.flag = "-lLLVMCodeGen",
    core.linker.flag = "-lLLVMCodeGenTypes",
    core.linker.flag = "-lLLVMCore",
    core.linker.flag = "-lLLVMCoroutines",
    core.linker.flag = "-lLLVMCoverage",
    core.linker.flag = "-lLLVMDebugInfoBTF",
    core.linker.flag = "-lLLVMDebugInfoCodeView",
    core.linker.flag = "-lLLVMDebuginfod",
    core.linker.flag = "-lLLVMDebugInfoDWARF",
    core.linker.flag = "-lLLVMDebugInfoDWARFLowLevel",
    core.linker.flag = "-lLLVMDebugInfoGSYM",
    core.linker.flag = "-lLLVMDebugInfoLogicalView",
    core.linker.flag = "-lLLVMDebugInfoMSF",
    core.linker.flag = "-lLLVMDebugInfoPDB",
    core.linker.flag = "-lLLVMDemangle",
    core.linker.flag = "-lLLVMDiff",
    core.linker.flag = "-lLLVMDlltoolDriver",
    core.linker.flag = "-lLLVMDWARFLinker",
    core.linker.flag = "-lLLVMDWARFLinkerClassic",
    core.linker.flag = "-lLLVMDWARFLinkerParallel",
    core.linker.flag = "-lLLVMDWP",
    core.linker.flag = "-lLLVMExecutionEngine",
    core.linker.flag = "-lLLVMExegesis",
    core.linker.flag = "-lLLVMExegesisAArch64",
    core.linker.flag = "-lLLVMExegesisMips",
    core.linker.flag = "-lLLVMExegesisPowerPC",
    core.linker.flag = "-lLLVMExegesisX86",
    core.linker.flag = "-lLLVMExtensions",
    core.linker.flag = "-lLLVMFileCheck",
    core.linker.flag = "-lLLVMFrontendAtomic",
    core.linker.flag = "-lLLVMFrontendDriver",
    core.linker.flag = "-lLLVMFrontendHLSL",
    core.linker.flag = "-lLLVMFrontendOffloading",
    core.linker.flag = "-lLLVMFrontendOpenACC",
    core.linker.flag = "-lLLVMFrontendOpenMP",
    core.linker.flag = "-lLLVMFuzzerCLI",
    core.linker.flag = "-lLLVMFuzzMutate",
    core.linker.flag = "-lLLVMGlobalISel",
    core.linker.flag = "-lLLVMHexagonAsmParser",
    core.linker.flag = "-lLLVMHexagonCodeGen",
    core.linker.flag = "-lLLVMHexagonDesc",
    core.linker.flag = "-lLLVMHexagonDisassembler",
    core.linker.flag = "-lLLVMHexagonInfo",
    core.linker.flag = "-lLLVMHipStdPar",
    core.linker.flag = "-lLLVMInstCombine",
    core.linker.flag = "-lLLVMInstrumentation",
    core.linker.flag = "-lLLVMInterfaceStub",
    core.linker.flag = "-lLLVMInterpreter",
    core.linker.flag = "-lLLVMipo",
    core.linker.flag = "-lLLVMIRPrinter",
    core.linker.flag = "-lLLVMIRReader",
    core.linker.flag = "-lLLVMJITLink",
    core.linker.flag = "-lLLVMLanaiAsmParser",
    core.linker.flag = "-lLLVMLanaiCodeGen",
    core.linker.flag = "-lLLVMLanaiDesc",
    core.linker.flag = "-lLLVMLanaiDisassembler",
    core.linker.flag = "-lLLVMLanaiInfo",
    core.linker.flag = "-lLLVMLibDriver",
    core.linker.flag = "-lLLVMLineEditor",
    core.linker.flag = "-lLLVMLinker",
    core.linker.flag = "-lLLVMLoongArchAsmParser",
    core.linker.flag = "-lLLVMLoongArchCodeGen",
    core.linker.flag = "-lLLVMLoongArchDesc",
    core.linker.flag = "-lLLVMLoongArchDisassembler",
    core.linker.flag = "-lLLVMLoongArchInfo",
    core.linker.flag = "-lLLVMLTO",
    core.linker.flag = "-lLLVMMC",
    core.linker.flag = "-lLLVMMCA",
    core.linker.flag = "-lLLVMMCDisassembler",
    core.linker.flag = "-lLLVMMCJIT",
    core.linker.flag = "-lLLVMMCParser",
    core.linker.flag = "-lLLVMMipsAsmParser",
    core.linker.flag = "-lLLVMMipsCodeGen",
    core.linker.flag = "-lLLVMMipsDesc",
    core.linker.flag = "-lLLVMMipsDisassembler",
    core.linker.flag = "-lLLVMMipsInfo",
    core.linker.flag = "-lLLVMMIRParser",
    core.linker.flag = "-lLLVMMSP430AsmParser",
    core.linker.flag = "-lLLVMMSP430CodeGen",
    core.linker.flag = "-lLLVMMSP430Desc",
    core.linker.flag = "-lLLVMMSP430Disassembler",
    core.linker.flag = "-lLLVMMSP430Info",
    core.linker.flag = "-lLLVMNVPTXCodeGen",
    core.linker.flag = "-lLLVMNVPTXDesc",
    core.linker.flag = "-lLLVMNVPTXInfo",
    core.linker.flag = "-lLLVMObjCARCOpts",
    core.linker.flag = "-lLLVMObjCopy",
    core.linker.flag = "-lLLVMObject",
    core.linker.flag = "-lLLVMObjectYAML",
    core.linker.flag = "-lLLVMOptDriver",
    core.linker.flag = "-lLLVMOption",
    core.linker.flag = "-lLLVMOrcDebugging",
    core.linker.flag = "-lLLVMOrcJIT",
    core.linker.flag = "-lLLVMOrcShared",
    core.linker.flag = "-lLLVMOrcTargetProcess",
    core.linker.flag = "-lLLVMPasses",
    core.linker.flag = "-lLLVMPowerPCAsmParser",
    core.linker.flag = "-lLLVMPowerPCCodeGen",
    core.linker.flag = "-lLLVMPowerPCDesc",
    core.linker.flag = "-lLLVMPowerPCDisassembler",
    core.linker.flag = "-lLLVMPowerPCInfo",
    core.linker.flag = "-lLLVMProfileData",
    core.linker.flag = "-lLLVMRemarks",
    core.linker.flag = "-lLLVMRISCVAsmParser",
    core.linker.flag = "-lLLVMRISCVCodeGen",
    core.linker.flag = "-lLLVMRISCVDesc",
    core.linker.flag = "-lLLVMRISCVDisassembler",
    core.linker.flag = "-lLLVMRISCVInfo",
    core.linker.flag = "-lLLVMRISCVTargetMCA",
    core.linker.flag = "-lLLVMRuntimeDyld",
    core.linker.flag = "-lLLVMSandboxIR",
    core.linker.flag = "-lLLVMScalarOpts",
    core.linker.flag = "-lLLVMSelectionDAG",
    core.linker.flag = "-lLLVMSparcAsmParser",
    core.linker.flag = "-lLLVMSparcCodeGen",
    core.linker.flag = "-lLLVMSparcDesc",
    core.linker.flag = "-lLLVMSparcDisassembler",
    core.linker.flag = "-lLLVMSparcInfo",
    core.linker.flag = "-lLLVMSPIRVAnalysis",
    core.linker.flag = "-lLLVMSPIRVCodeGen",
    core.linker.flag = "-lLLVMSPIRVDesc",
    core.linker.flag = "-lLLVMSPIRVInfo",
    core.linker.flag = "-lLLVMSupport",
    core.linker.flag = "-lLLVMSymbolize",
    core.linker.flag = "-lLLVMSystemZAsmParser",
    core.linker.flag = "-lLLVMSystemZCodeGen",
    core.linker.flag = "-lLLVMSystemZDesc",
    core.linker.flag = "-lLLVMSystemZDisassembler",
    core.linker.flag = "-lLLVMSystemZInfo",
    core.linker.flag = "-lLLVMTableGen",
    core.linker.flag = "-lLLVMTableGenBasic",
    core.linker.flag = "-lLLVMTableGenCommon",
    core.linker.flag = "-lLLVMTarget",
    core.linker.flag = "-lLLVMTargetParser",
    core.linker.flag = "-lLLVMTelemetry",
    core.linker.flag = "-lLLVMTextAPI",
    core.linker.flag = "-lLLVMTextAPIBinaryReader",
    core.linker.flag = "-lLLVMTransformUtils",
    core.linker.flag = "-lLLVMVEAsmParser",
    core.linker.flag = "-lLLVMVECodeGen",
    core.linker.flag = "-lLLVMVectorize",
    core.linker.flag = "-lLLVMVEDesc",
    core.linker.flag = "-lLLVMVEDisassembler",
    core.linker.flag = "-lLLVMVEInfo",
    core.linker.flag = "-lLLVMWebAssemblyAsmParser",
    core.linker.flag = "-lLLVMWebAssemblyCodeGen",
    core.linker.flag = "-lLLVMWebAssemblyDesc",
    core.linker.flag = "-lLLVMWebAssemblyDisassembler",
    core.linker.flag = "-lLLVMWebAssemblyInfo",
    core.linker.flag = "-lLLVMWebAssemblyUtils",
    core.linker.flag = "-lLLVMWindowsDriver",
    core.linker.flag = "-lLLVMWindowsManifest",
    core.linker.flag = "-lLLVMX86AsmParser",
    core.linker.flag = "-lLLVMX86CodeGen",
    core.linker.flag = "-lLLVMX86Desc",
    core.linker.flag = "-lLLVMX86Disassembler",
    core.linker.flag = "-lLLVMX86Info",
    core.linker.flag = "-lLLVMX86TargetMCA",
    core.linker.flag = "-lLLVMXCoreCodeGen",
    core.linker.flag = "-lLLVMXCoreDesc",
    core.linker.flag = "-lLLVMXCoreDisassembler",
    core.linker.flag = "-lLLVMXCoreInfo",
    core.linker.flag = "-lLLVMXRay",
    core.linker.flag = "-lstdc++",
    core.linker.flag = "-pthread",
    // Wrapper around target macro definitions
    core.linker.additionalSource = "target-wrapper.c"
]
