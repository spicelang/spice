f<int> main() {
    assert 1 != 1;
    printf("Unreachable");
}