public type IScope interface {

}