type T dyn;

f<T> test() {
    return 1;
}

f<int> main() {
    test();
}