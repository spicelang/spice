type TokenType enum {
    IDENTIFIER,
    DOT = 12,
    COMMA,
    SIZEOF = 0,
    WS
}

f<int> main() {
    printf("%d\n", TokenType::DOT);
    printf("%d\n", TokenType::COMMA);
    printf("%d\n", TokenType::IDENTIFIER);
    printf("%d\n", TokenType::WS);
    printf("%d\n", TokenType::SIZEOF);
}