import "../../src-bootstrap/reader/reader";

f<int> main() {
    Reader reader = Reader("./test.spice");
}