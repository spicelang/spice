unsigned short unsignedShort = -10;
const signed int test = 6s;

f<int> main() {
    printf("Int: %d", test);
}