// Converts an int to a double
f<double> toDouble(int input) {
    // ToDo: Implement
    return 0.0;
}

// Converts an int to a byte
f<type> toDouble(int input) {
    // ToDo: Implement
    return 0 + input;
}

// Converts an int to a char
f<char> ToByte(int input) {
    // ToDo: Implement
    result = 0 + input;
}

// Converts an int to a char
f<char> ToChar(int input) {
    // ToDo: Implement
    return 0 + input;
}

// Converts an int to a string
f<string> toString(int input) {
    // ToDo: Implement (See https://github.com/golang/go/blob/master/src/strconv/itoa.go)
    return "";
}

// Converts an int to a boolean
f<bool> toBool(int input) {
    return input >= 1;
}