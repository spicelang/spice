import "std/type/result";

// Add generic type definitions
type K dyn;
type V dyn;

// Enums
type NodeColor enum { RED, BLACK }

/**
 * Node of a Red-Black Tree
 */
type Node<K, V> struct {
    K key
    V value
    NodeColor color
    heap Node<K, V>* parent
    heap Node<K, V>* childLeft
    heap Node<K, V>* childRight
}

inline f<bool> Node.isRoot() {
    return this.parent == nil<heap Node<K, V>*>;
}

/**
 * A Red-Black Tree is a self-balancing search tree, which is used e.g. in the implementation of maps.
 *
 * Time complexity:
 * Insert: O(log n)
 * Delete: O(log n)
 * Lookup: O(log n)
 */
public type RedBlackTree<K, V> struct {
    heap Node<K, V>* rootNode
}

public p RedBlackTree.ctor() {
    this.rootNode = nil<heap Node<K, V>*>;
}

p RedBlackTree.rotateLeft(heap Node<K, V>* x) {
    heap Node<K, V>* y = x.childRight;
    x.childRight = y.childLeft;
    if y.childLeft != nil<heap Node<K, V>*> {
        y.childLeft.parent = x;
    }
    y.parent = x.parent;
    if x.parent == nil<heap Node<K, V>*> {
        this.rootNode = y;
    } else if x == x.parent.childLeft {
        x.parent.childLeft = y;
    } else {
        x.parent.childRight = y;
    }
    y.childLeft = x;
    x.parent = y;
}

p RedBlackTree.rotateRight(heap Node<K, V>* y) {
    heap Node<K, V>* x = y.childLeft;
    y.childLeft = x.childRight;
    if x.childRight != nil<heap Node<K, V>*> {
        x.childRight.parent = y;
    }
    x.parent = y.parent;
    if y.parent == nil<heap Node<K, V>*> {
        this.rootNode = x;
    } else if y == y.parent.childRight {
        y.parent.childRight = x;
    } else {
        y.parent.childLeft = x;
    }
    x.childRight = y;
    y.parent = x;
}

p RedBlackTree.insertFixup(heap Node<K, V>* z) {
    while z.parent != nil<heap Node<K, V>*> && z.parent.color == NodeColor::RED {
        if z.parent == z.parent.parent.childLeft {
            heap Node<K, V>* y = z.parent.parent.childRight;
            if y != nil<heap Node<K, V>*> && y.color == NodeColor::RED {
                z.parent.color = NodeColor::BLACK;
                y.color = NodeColor::BLACK;
                z.parent.parent.color = NodeColor::RED;
                z = z.parent.parent;
            } else {
                if z == z.parent.childRight {
                    z = z.parent;
                    this.rotateLeft(z);
                }
                z.parent.color = NodeColor::BLACK;
                z.parent.parent.color = NodeColor::RED;
                this.rotateRight(z.parent.parent);
            }
        } else {
            heap Node<K, V>* y = z.parent.parent.childLeft;
            if y != nil<heap Node<K, V>*> && y.color == NodeColor::RED {
                z.parent.color = NodeColor::BLACK;
                y.color = NodeColor::BLACK;
                z.parent.parent.color = NodeColor::RED;
                z = z.parent.parent;
            } else {
                if z == z.parent.childLeft {
                    z = z.parent;
                    this.rotateRight(z);
                }
                z.parent.color = NodeColor::BLACK;
                z.parent.parent.color = NodeColor::RED;
                this.rotateLeft(z.parent.parent);
            }
        }
    }
    this.rootNode.color = NodeColor::BLACK;
}

p RedBlackTree.transplant(heap Node<K, V>* u, heap Node<K, V>* v) {
    if u.parent == nil<heap Node<K, V>*> {
        this.rootNode = v;
    } else if u == u.parent.childLeft {
        u.parent.childLeft = v;
    } else {
        u.parent.childRight = v;
    }
    if v != nil<heap Node<K, V>*> {
        v.parent = u.parent;
    }
}

p RedBlackTree.deleteFixup(heap Node<K, V>* x) {
    while x != this.rootNode && (x == nil<Node<K, V>*> || x.color == NodeColor::BLACK) {
        if x == x.parent.childLeft {
            Node<K, V>* w = x.parent.childRight;
            if w != nil<Node<K, V>*> && w.color == NodeColor::RED {
                w.color = NodeColor::BLACK;
                x.parent.color = NodeColor::RED;
                this.rotateLeft(x.parent);
                w = x.parent.childRight;
            }
            if (w.childLeft == nil<Node<K, V>*> || w.childLeft.color == NodeColor::BLACK) && (w.childRight == nil<Node<K, V>*> || w.childRight.color == NodeColor::BLACK) {
                w.color = NodeColor::RED;
                x = x.parent;
            } else {
                if w.childRight == nil<Node<K, V>*> || w.childRight.color == NodeColor::BLACK {
                    if w.childLeft != nil<Node<K, V>*> {
                        w.childLeft.color = NodeColor::BLACK;
                    }
                    w.color = NodeColor::RED;
                    this.rotateRight(w);
                    w = x.parent.childRight;
                }
                w.color = x.parent.color;
                x.parent.color = NodeColor::BLACK;
                if w.childRight != nil<Node<K, V>*> {
                    w.childRight.color = NodeColor::BLACK;
                }
                this.rotateLeft(x.parent);
                x = this.rootNode;
            }
        } else {
            Node<K, V>* w = x.parent.childLeft;
            if w != nil<Node<K, V>*> && w.color == NodeColor::RED {
                w.color = NodeColor::BLACK;
                x.parent.color = NodeColor::RED;
                this.rotateRight(x.parent);
                w = x.parent.childLeft;
            }
            if (w.childRight == nil<Node<K, V>*> || w.childRight.color == NodeColor::BLACK) && (w.childLeft == nil<Node<K, V>*> || w.childLeft.color == NodeColor::BLACK) {
                w.color = NodeColor::RED;
                x = x.parent;
            } else {
                if w.childLeft == nil<Node<K, V>*> || w.childLeft.color == NodeColor::BLACK {
                    if w.childRight != nil<Node<K, V>*> {
                        w.childRight.color = NodeColor::BLACK;
                    }
                    w.color = NodeColor::RED;
                    this.rotateLeft(w);
                    w = x.parent.childLeft;
                }
                w.color = x.parent.color;
                x.parent.color = NodeColor::BLACK;
                if w.childLeft != nil<Node<K, V>*> {
                    w.childLeft.color = NodeColor::BLACK;
                }
                this.rotateRight(x.parent);
                x = this.rootNode;
            }
        }
    }
    if x != nil<Node<K, V>*> {
        x.color = NodeColor::BLACK;
    }
}

public p RedBlackTree.insert(const K& key, const V& value) {
    heap Node<K, V>* newNode = sNew<Node<K, V>>(Node<K, V>{
        key,
        value,
        NodeColor::RED,
        nil<heap Node<K, V>*>,
        nil<heap Node<K, V>*>,
        nil<heap Node<K, V>*>
    });
    heap Node<K, V>* y = nil<heap Node<K, V>*>;
    heap Node<K, V>* x = this.rootNode;
    while x != nil<heap Node<K, V>*> {
        y = x;
        if newNode.key < x.key {
            x = x.childLeft;
        } else {
            x = x.childRight;
        }
    }
    newNode.parent = y;
    if y == nil<heap Node<K, V>*> {
        this.rootNode = newNode;
    } else if newNode.key < y.key {
        y.childLeft = newNode;
    } else {
        y.childRight = newNode;
    }
    this.insertFixup(newNode);
}

public p RedBlackTree.remove(const K& key) {
    heap Node<K, V>* z = this.search(key);
    if z == nil<heap Node<K, V>*> {
        return;
    }
    heap Node<K, V>* y = z;
    heap Node<K, V>* x;
    NodeColor yOriginalColor = y.color;
    if z.childLeft == nil<heap Node<K, V>*> {
        x = z.childRight;
        this.transplant(z, z.childRight);
    } else if z.childRight == nil<heap Node<K, V>*> {
        x = z.childLeft;
        this.transplant(z, z.childLeft);
    } else {
        y = this.minimum(z.childRight);
        yOriginalColor = y.color;
        x = y.childRight;
        if y.parent == z {
            x.parent = y;
        } else {
            this.transplant(y, y.childRight);
            y.childRight = z.childRight;
            y.childRight.parent = y;
        }
        this.transplant(z, y);
        y.childLeft = z.childLeft;
        y.childLeft.parent = y;
        y.color = z.color;
    }
    sDelete(z);
    if yOriginalColor == NodeColor::BLACK {
        deleteFixup(x);
    }
}

public f<V&> RedBlackTree.find(const K& key) {
    return this.search(key).value;
}

public f<Result<V&>> RedBlackTree.findSafe(const K& key) {
    heap Node<K, V>* node = this.search(key);
    return node != nil<heap Node<K, V>*> ? ok(node.value) : err(Error("The provided key was not found"));
}

f<heap Node<K, V>*> RedBlackTree.search(const K& key) {
    heap Node<K, V>* currentNode = this.rootNode;
    while currentNode != nil<heap Node<K, V>*> {
        if key == currentNode.key {
            return currentNode;
        } else if key < currentNode.key {
            currentNode = currentNode.childLeft;
        } else {
            currentNode = currentNode.childRight;
        }
    }
    return nil<heap Node<K, V>*>;
}

public f<heap Node<K, V>*> RedBlackTree.minimum(heap Node<K, V>* x) {
    while x.childLeft != nil<heap Node<K, V>*> {
        x = x.childLeft;
    }
    return x;
}