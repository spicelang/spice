f<int> main() {
    double doubleVar = 1.34;
    doubleVar.test = 1;
}