public const unsigned int ANONYMOUS = 0;