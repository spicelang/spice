import "std/time/timer";

f<int> fibo(int n) {
    if n <= 1 { return n; }
    return fibo(n - 1) + fibo(n - 2);
}

f<int> main() {
    Timer t = Timer();
    t.start();
    printf("Output: %d\n", fibo(45));
    t.stop();
    printf("Elapsed time: %d\n", t.getDurationInMicros());
    printf("Elapsed time: %d\n", t.getDurationInMillis());
    printf("Elapsed time: %f\n", t.getDurationInSeconds());
    printf("Elapsed time: %f\n", t.getDurationInMinutes());
}