import "std/data/hash-table";
import "std/iterator/iterable";
import "std/iterator/iterator";
import "std/data/pair";

// Add generic type definitions
type K dyn;
type V dyn;

/**
 * An unordered map in Spice is a commonly used data structure, which can be used to represent a list of key value pairs.
 *
 * Time complexity:
 * Insert: O(1) (average case), O(n) (worst case)
 * Delete: O(1) (average case), O(n) (worst case)
 * Lookup: O(1) (average case), O(n) (worst case)
 */
public type UnorderedMap<K, V> struct : IIterable<Pair<K, V>> {
    HashTable<K, V> hashTable
}

public p UnorderedMap.ctor(unsigned long bucketCount = 100l) {
    this.hashTable = HashTable<K, V>(bucketCount);
}

/**
 * Insert a key-value pair into the map
 * If the key already exists, the value is updated.
 *
 * @param key The key to insert
 * @param value The value to insert
 */
public p UnorderedMap.upsert(const K& key, const V& value) {
    this.hashTable.upsert(key, value);
}

/**
 * Retrieve the value associated with the given key.
 * If the key is not found, panic.
 *
 * @param key The key to look up
 * @return The value associated with the key
 */
public f<V&> UnorderedMap.get(const K& key) {
    return this.hashTable.get(key);
}

/**
 * Retrieve the value associated with the given key.
 * If the key is not found, panic.
 *
 * @param key The key to look up
 * @return The value associated with the key
 */
public f<V&> operator[]<K, V>(UnorderedMap<K, V>& map, const K& key) {
    return map.get(key);
}

/**
 * Retrieve the value associated with the given key as Result<V>.
 * If the key is not found, the result contains an error.
 *
 * @param key The key to look up
 * @return Result<V>, containing the value associated with the key or an error if the key is not found
 */
public f<Result<V>> UnorderedMap.getSafe(const K& key) {
    return this.hashTable.getSafe(key);
}

/**
 * Check if the map contains the given key.
 *
 * @param key The key to check for
 * @return True if the key is found, false otherwise
 */
public p UnorderedMap.remove(const K& key) {
    this.hashTable.remove(key);
}

/**
 * Check if the map contains the given key.
 *
 * @param key The key to check for
 * @return True if the key is found, false otherwise
 */
public f<bool> UnorderedMap.contains(const K& key) {
    return this.hashTable.contains(key);
}

/**
 * Get the size of the unordered map.
 *
 * @return The number of key-value pairs in the map
 */
public f<unsigned long> UnorderedMap.getSize() {
    return this.hashTable.getSize();
}

/**
 * Check if the unordered map is empty.
 *
 * @return True if empty, false otherwise
 */
public f<bool> UnorderedMap.isEmpty() {
    return this.hashTable.isEmpty();
}

/**
 * Clear the unordered map, removing all key-value pairs.
 */
public p UnorderedMap.clear() {
    this.hashTable.clear();
}

/**
 * Iterator to iterate over an unordered map data structure
 */
public type UnorderedMapIterator<K, V> struct : IIterator<Pair<const K&, V&>> {
    HashTableIterator<K, V> htIterator
}

public p UnorderedMapIterator.ctor<K, V>(UnorderedMap<K, V>& unorderedMap) {
    this.htIterator = unorderedMap.hashTable.getIterator();
}
/**
 * Returns the current key-value pair of the unordered map
 *
 * @return Current key/value pair
 */
public inline f<Pair<const K&, V&>&> UnorderedMapIterator.get() {
    return this.htIterator.get();
}

/**
 * Returns the current index and the current item of the unordered map
 *
 * @return Pair of current index and current key/value pair
 */
public inline f<Pair<unsigned long, Pair<const K&, V&>&>> UnorderedMapIterator.getIdx() {
    return this.htIterator.getIdx();
}

/**
 * Check if the iterator is valid
 *
 * @return true or false
 */
public inline f<bool> UnorderedMapIterator.isValid() {
    return this.htIterator.isValid();
}

/**
 * Moves the cursor to the next key/value pair
 */
public inline p UnorderedMapIterator.next() {
    this.htIterator.next();
}

/**
 * Advances the cursor by one
 *
 * @param it UnorderedMapIterator
 */
public inline p operator++<K, V>(UnorderedMapIterator<K, V>& it) {
    this.htIterator.next();
}

/**
 * Retrieve a forward iterator for the unordered map
 */
public f<UnorderedMapIterator<K, V>> UnorderedMap.getIterator() {
    return UnorderedMapIterator<K, V>(*this);
}
