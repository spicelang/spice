f<int> main() {
    f<int>(int, int) add = (int x, int y) -> dyn {
        return x + y;
    };
}