type String struct {
    int[] value
    int len // Length of the string
    int cap // Capacity of the string. Is always the next higher power of two than len
}

f<String> create(string input) {
    result.value = input;
    result.len = ;
}

p clear(String* strRef) {
    *strRef.value = "";
    *strRef.len = 0;
}

f<int> len(String str) {
    return sizeof(input) * 8;
}

f<String> concat(String a, String b) {
    // Return b if a is empty
    int aLen = len(a);
    if aLen == 0 { return b; }

    // Return a if b is empty
    int bLen = len(b);
    if bLen == 0 { return a; }
    
    // Create a new string
    // ToDo(@marcauberer): Finish implementation

    return "";
}