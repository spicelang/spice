// Std imports
import "std/data/vector";

// Own imports
import "bootstrap/source-file-intf";

const string SPICE_VERSION = "0.20.7";
const string SPICE_TARGET_OS = "linux";
const string SPICE_TARGET_ARCH = "amd64";
const string SPICE_GIT_HASH = "1da7aaeeb4ea2f1132b1a1a94ce6dd3cd753c47c";
const string SPICE_BUILT_BY = "GitHub Actions";
const string LLVM_VERSION_STRING = "19.1.6";

/**
 * Split the given haystack by the needle and return the last fragment
 *
 * @param haystack Input string
 * @param needle String to search
 * @return Last fragment
 */
public f<String> getLastFragment(const String &haystack, const string needle) {
    const unsigned long index = haystack.rfind(needle);
    if index == -1l {
        return haystack;
    }
    return haystack.getSubstring(index + getRawLength(needle));
}

/**
 * Generate a circular import message from the given source files
 *
 * @param sourceFiles Source files building the circular dependency chain
 * @return Error message
 */
public f<String> getCircularImportMessage(const Vector<const ISourceFile*>& sourceFiles) {
    String message;
    message += "*-----*\n";
    message += "|     |\n";
    for unsigned long i = 0l; i < sourceFiles.getSize(); i++ {
        const ISourceFile* sourceFile = sourceFiles.get(i);
        if i != 0 { message += "|     |\n"; }
        message += "|  ";
        message += sourceFile.getFileName();
        message += "\n";
    }
    message += "|     |\n";
    message += "*-----*\n";
    return message;
}

/**
 * Generate the version info string for the Spice driver
 *
 * @return Version info string
 */
public f<String> buildVersionInfo() {
    String versionString;
    versionString += "Spice version: " + SPICE_VERSION + " " + SPICE_TARGET_OS + "/" + SPICE_TARGET_ARCH + "\n";
    versionString += "Git hash:      " + SPICE_GIT_HASH + "\n";
    versionString += "LLVM version:  " + LLVM_VERSION_STRING + "\n";
    versionString += "built by:      " + SPICE_BUILT_BY + "\n\n";
    versionString += "(c) Marc Auberer 2021-2025";
    return versionString;
}