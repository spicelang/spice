f<int> main() {
    int i = 0;
    while i < 10 {
        i += 1;
        printf("i is now at: %d\n", i);
        if i > 5 {
            continue;
        }
        printf("test");
    }
}