import "std/runtime/string_rt" as _rt_str;

f<int> main() {
    _rt_str::String s = _rt_str::String('H');
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.append("ello");
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d", s.getCapacity());
}