public type SuperType enum {
    TY_INVALID,
    TY_UNRESOLVED,
    TY_DOUBLE,
    TY_INT,
    TY_SHORT,
    TY_LONG,
    TY_BYTE,
    TY_CHAR,
    TY_STRING, // Alias for 'const char*'
    TY_BOOL,
    TY_STRUCT,
    TY_INTERFACE,
    TY_ENUM,
    TY_GENERIC,
    TY_ALIAS,
    TY_DYN,
    TY_PTR,
    TY_REF,
    TY_ARRAY,
    TY_FUNCTION,
    TY_PROCEDURE,
    TY_IMPORT
}