p test() {
    printf("Test called.");
    return "Invalid return value";
}

f<int> main() {
    test();
}