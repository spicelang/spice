public p test() {
    printf("Hello World");
}