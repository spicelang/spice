type Struct struct {
    const int& ref
}

f<int> main() {
    int i = 123;
    Struct str = Struct { 123 };
    printf("Field value: %d", str.ref);
}