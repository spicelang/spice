p testProc(string arg0, bool arg1 = false, int arg2) {
    printf("Test");
}

f<int> main() {
    testProc("test", true);
}