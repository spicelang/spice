#![core.linker.additionalSource = "non-existing.c"]

f<int> main() {
    testFunction();
}