type T string|const char*;

p foo<T>(T str) {}

f<int> main() {
    foo(cast<const char*>("hello"));
    foo("world");
}