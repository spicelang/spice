import "std/io/cli-parser";

type CliOptions struct {
    string greetName = ""
}

p callback(bool& value) {
    printf("Callback called with value %d\n", value);
}

f<int> main(int argc, string[] argv) {
    CliParser parser = CliParser("Test Program", "This is a simple test program");
    parser.setVersion("v0.1.0");
    parser.setFooter("Copyright (c) Marc Auberer 2021-2023");

    CliOptions options;
    CliSubcommand& greet = parser.addSubcommand("greet", "Greet someone");
    greet.addOption("--name", options.greetName, "Name of the person to greet");

    parser.parse(argc, argv);

    // Greet persion if requested
    if options.greetName != "" {
        printf("Hello %s!\n", options.greetName);
    }
}