public type TestStruct struct {

}