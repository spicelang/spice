f<int> main() {}