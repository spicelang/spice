public const int SIZE = 8;
public const int MIN_VALUE = 0;
public const int MAX_VALUE = 255;

// Converts a char to a double
public f<double> toDouble(char input) {
    return 0.0 + (int) input;
}

// Converts a char to an int
public f<int> toInt(char input) {
    return (int) input;
}

// Converts a char to a short
public f<short> toShort(char input) {
    return (short) ((int) input);
}

// Converts a char to a long
public f<long> toLong(char input) {
    return (long) ((int) input);
}

// Converts a char to a byte
public f<byte> toByte(char input) {
    result = (byte) input;
}

// Converts a char to a string
public f<String> toString(char input) {
    result = String();
    result += input;
}

// Converts a char to a bool
public f<bool> toBool(char input) {
    return input == '1';
}