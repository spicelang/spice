f<int> main() {
    printf("%f", true);
}