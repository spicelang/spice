f<int> main() {
    if ("test" || false) {
        printf("Hello World!");
    }
    if (true && 6) {
        printf("Hello World!");
    }
}