f<bool> cond1() {
    printf("cond1");
    return true;
}

f<bool> cond2() {
    printf("cond2");
    return true;
}

f<bool> cond3() {
    printf("cond3");
    return true;
}

f<int> main() {
    if cond1() && cond2() && cond3() {
        printf("true");
        return 0;
    }
    printf("false");
}