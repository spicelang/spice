import "std/iterator/iterator";
import "std/data/pair";

// Generic type definitions
type I dyn;
type Numeric int|long|short;

/**
 * An ArrayIterator in Spice can be used to iterate over an arbitrary array
 */
public type ArrayIterator<I> struct : IIterator<I> {
    I* array
    unsigned long size
    unsigned long cursor = 0l
}

public p ArrayIterator.ctor(I[] array, unsigned long size) {
    this.array = array;
    this.size = size;
}

/**
 * Returns the current item of the array
 *
 * @return Reference to the current item
 */
public inline f<I&> ArrayIterator.get() {
    unsafe {
        return this.array[this.cursor];
    }
}

public inline f<Pair<unsigned long, I&>> ArrayIterator.getIdx() {
    unsafe {
        return Pair<unsigned long, I&>(this.cursor, this.array[this.cursor]);
    }
}

/**
 * Check if the iterator is valid
 *
 * @return true or false
 */
public inline const f<bool> ArrayIterator.isValid() {
    return this.cursor < this.size;
}

/**
 * Returns the current item of the array and moves the cursor to the next one
 */
public inline p ArrayIterator.next() {
    if !this.isValid() { panic(Error("Calling next() on invalid iterator")); }
    this.cursor++;
}

/**
 * Advances the cursor by one
 *
 * @param it ArrayIterator
 */
public inline p operator++<I>(ArrayIterator<I>& it) {
    if it.cursor >= it.size - 1l { panic(Error("Iterator out of bounds")); }
    it.cursor++;
}

/**
 * Move the cursor back by one
 *
 * @param it ArrayIterator
 */
public inline p operator--<I>(ArrayIterator<I>& it) {
    if it.cursor <= 0l { panic(Error("Iterator out of bounds")); }
    it.cursor--;
}

/**
 * Advances the cursor by the given offset
 *
 * @param it ArrayIterator
 * @param offset Offset
 */
public inline p operator+=<I, Numeric>(ArrayIterator<I>& it, Numeric offset) {
    if it.cursor + offset >= it.size || it.cursor + offset < 0l { panic(Error("Iterator out of bounds")); }
    it.cursor += offset;
}

/**
 * Move the cursor back by the given offset
 *
 * @param it ArrayIterator
 * @param offset Offset
 */
public inline p operator-=<I, Numeric>(ArrayIterator<I>& it, Numeric offset) {
    if it.cursor - offset >= it.size || it.cursor - offset < 0l { panic(Error("Iterator out of bounds")); }
    it.cursor -= offset;
}

/**
 * Convenience wrapper for creating a simple array iterator
 */
public inline f<ArrayIterator<I>> iterate<I>(I[] array, unsigned long size) {
    return ArrayIterator<I>(array, size);
}