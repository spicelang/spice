f<int> main() {
    string test = "Tested";
    printf("%s\n", test.getRaw());
    printf("%d\n", test.getLength());
    printf("%d\n", test.getCapacity());
}

/*f<int> main() {
    int v1 = 10;
    int v2 = v1;
    printf("v1: %d, v2: %d\n", v1, v2);
    v2++;
    printf("v1: %d, v2: %d\n", v1, v2);

    unsigned long startIndex = 10l;
    for unsigned long charIndex = startIndex; charIndex < 20l; charIndex++ {
        printf("Char index: %d, start index: %d\n", charIndex, startIndex);
    }
}*/

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

/*public f<bool> src(bool x, bool y) {
    return ((x ? 1 : 4) & (y ? 1 : 4)) == 0;
}

public f<int> tgt(int x, int y) {
    return x ^ y;
}

f<int> main() {
    printf("Result: %d, %d", src(false, true), tgt(0, 1));
}*/