// Std imports

// Own imports

public type ISourceFile interface {
    public f<unsigned long> getLineCount();
    public f<string> getFileName();
}