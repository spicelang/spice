f<int> main() {
    do {
        printf("Test");
    } while(5.6);
}