import "test2" as s1;

f<int> main() {
    s1.test();
}

f<double> getDouble() {
    return 4.3;
}