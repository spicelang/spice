/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec.Vector<pair.Pair<int, string>> pairVector = vec.Vector<pair.Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair.Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

/*const unsigned int vertexCount = 9;

f<int> main() {
    int[vertexCount][vertexCount] graph = {
        { 0, 4, 0, 0, 0, 0, 0, 8, 0 },
        { 4, 0, 8, 0, 0, 0, 0, 11, 0 },
        { 0, 8, 0, 7, 0, 4, 0, 0, 2 },
        { 0, 0, 7, 0, 9, 14, 0, 0, 0 },
        { 0, 0, 0, 9, 0, 10, 0, 0, 0 },
        { 0, 0, 4, 14, 10, 0, 2, 0, 0 },
        { 0, 0, 0, 0, 0, 2, 0, 1, 6 },
        { 8, 11, 0, 0, 0, 0, 1, 0, 7 },
        { 0, 0, 2, 0, 0, 0, 6, 7, 0 }
    };

    printf("Test: %d, %d\n", graph[1][7], sizeof(graph));
}*/

/*f<int> main() {
    printf("Array1:\n");
    short arraySize1 = 4s;
    int[arraySize1] array1 = {1, 2, 3};
    array1[3] = 0;
    foreach dyn item : array1 {
        printf("Item: %d\n", item);
    }

    printf("Array2:\n");
    long arraySize2 = 2l;
    string[arraySize2] array2;
    array2[0] = "Hello";
    array2[1] = "world";
    foreach dyn item : array2 {
        printf("Item: %s\n", item);
    }

    printf("Array3:\n");
    int arraySize3 = 3;
    int[arraySize3] array3 = {1, arraySize3, arraySize3};
    foreach dyn item : array3 {
        printf("Item: %d\n", item);
    }

    printf("Array4:\n");
    int arraySize4 = 3;
    int[arraySize4] array4;
    array4 = {1, arraySize4, arraySize4};
    foreach dyn item : array4 {
        printf("Item: %d\n", item);
    }
}*/

int count = -5;

f<int> main() {
    int[count] items;
    /*items[0] = 1;
    items[1] = 2;
    items[2] = 3;
    items[3] = 4;
    items[4] = 5;*/
    foreach int i : items {
        printf("%d\n", i);
    }
}