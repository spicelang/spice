// Converts a string to a double
public f<double> toDouble(string input) {
    // ToDo: implement
    return 0.0;
}

// Converts a string to an int
public f<int> toInt(string input) {
    if input == "" {
        return 0;
    }

    bool neg = false;
    

    // ToDo: implement the rest
    return 0;
}

// Converts a string to a short
public f<short> toShort(string input) {
    if input == "" {
        return (short) 0;
    }

    bool neg = false;
    

    // ToDo: implement the rest
    return (short) 0;
}

// Converts a string to a long
public f<long> toLong(string input) {
    if input == "" {
        return (long) 0;
    }

    bool neg = false;
    

    // ToDo: implement the rest
    return (long) 0;
}

// Converts a string to a byte
public f<byte> toByte(string input) {
    if input == "" {
        return (byte) 0;
    }

    bool neg = false;
    

    // ToDo: implement the rest
    return (byte) 0;
}

// Converts a string to a char
public f<char> toChar(string input) {
    // ToDo: Implement
    return '0';
}

// Converts a string to a bool
public f<bool> toBool(string input) {
    return input == "true";
}

// Returns the length of a string
public f<long> getRawLength(string input) {
    result = 0l;
    while input[result] != '\0' {
        result++;
    }
}

// Returns the equality of two strings
public f<bool> isRawEqual(string lhs, string rhs) {
    unsigned long lhsLength = getRawLength(lhs);
    unsigned long rhsLength = getRawLength(rhs);
    // Return false immediately if length does not match
    if lhsLength != rhsLength { return false; }
    // Compare chars
    for int i = 0; i < lhsLength; i++ {
        if lhs[i] != rhs[i] {
            return false;
        }
    }
    return true;
}
