type Vector struct {
    int i
}