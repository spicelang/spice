// Std imports
import "std/os/os";

// Own imports
import "./source-file";
import "./driver";
import "./global/global-resource-manager";

/**
 * Compile main source file. All files, that are included by the main source file will be resolved recursively.
 *
 * @param cliOptions Command line options
 * @return Successful or not
 */
f<bool> compileProject(const CliOptions& cliOptions) {
    // Instantiate GlobalResourceManager
    dyn resourceManager = GlobalResourceManager(options);

    // Create source file instance for main source file
    SourceFile* mainSourceFile = resourceManager.createSourceFile(nullptr, MAIN_FILE_NAME, cliOptions.mainFile, false);

    // Run compile pipeline for main source file. All dependent source files are triggered by their parents
    mainSourceFile.runFrontEnd();
    mainSourceFile.runMiddleEnd();
    mainSourceFile.runBackEnd();

    // Link the target executable (link object files to executable)
    resourceManager.linker.prepare();
    resourceManager.linker.link();

    // Print compiler warnings
    mainSourceFile.collectAndPrintWarnings();

    // Print compiler warnings
    mainSourceFile.collectAndPrintWarnings();

    return true;
}

/**
 * Entry point to the Spice compiler
 *
 * @param argc Argument count
 * @param argv Argument vector
 * @return Return code
 */
f<int> main(int argc, string[] argv) {
    // Initialize command line parser
    Driver driver;
    driver.create();
    const int exitCode = driver.parse(argc, argv);
    if exitCode != EXIT_SUCCESS {
        return exitCode;
    }

    // Cancel here if we do not have to compile
    if !driver.shouldCompile {
        return EXIT_SUCCESS;
    }

    driver.enrich(); // Prepare the cli options

    // Kick off the compiling process
    if !compileProject(driver.cliOptions) {
        return EXIT_FAILURE;
    }

    // Execute
    if driver.cliOptions.execute {
        driver.runBinary();
    }

    return EXIT_SUCCESS;
}