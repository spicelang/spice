type TLhs dyn;
type TRhs dyn;

// ------------------------------------------ += ------------------------------------------

p plusEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs += rhs;
    assert lhs == expectedResult;
}

p plusEqualTestInnerUnsafe<TRhs>(int* lhs, const TRhs rhs, const int* expectedResult) {
    unsafe {
        lhs += rhs;
    }
    assert lhs == expectedResult;
}

p plusEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    plusEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    plusEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    plusEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    plusEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p plusEqualTest() {
    // Lhs is double
    plusEqualTestOuter<double, double>(1.234, 98.7654, 99.9994, -99.9994, 97.5314, -97.5314);
    // Lhs is int
    plusEqualTestOuter<int, int>(78, 674, 752, -752, 596, -596);
    plusEqualTestOuter<int, short>(78, 7s, 85, -85, -71, 71);
    plusEqualTestOuter<int, long>(78, 2384723l, 2384801, -2384801, 2384645, -2384645);
    // Lhs is short
    plusEqualTestOuter<short, int>(78s, 674, 752s, -752s, 596s, -596s);
    plusEqualTestOuter<short, short>(78s, 7s, 85s, -85s, -71s, 71s);
    plusEqualTestOuter<short, long>(78s, 2384723l, 25505s, -25505s, 25349s, -25349s);
    // Lhs is long
    plusEqualTestOuter<long, int>(78l, 674, 752l, -752l, 596l, -596l);
    plusEqualTestOuter<long, short>(78l, 7s, 85l, -85l, -71l, 71l);
    plusEqualTestOuter<long, long>(78l, 2384723l, 2384801l, -2384801l, 2384645l, -2384645l);
    // Lhs is char
    plusEqualTestInner<char, int>('A', 5, 'F');
    plusEqualTestInner<char, int>('A', -5, '<');
    // Lhs is ptr
    int[5] input = [0, 0, 0, 0, 0];
    plusEqualTestInnerUnsafe(&input[2], 2, &input[4]);
    plusEqualTestInnerUnsafe(&input[2], -2, &input[0]);
    plusEqualTestInnerUnsafe(&input[2], 2s, &input[4]);
    plusEqualTestInnerUnsafe(&input[2], -2s, &input[0]);
    plusEqualTestInnerUnsafe(&input[2], 2l, &input[4]);
    plusEqualTestInnerUnsafe(&input[2], -2l, &input[0]);
}

// ------------------------------------------ -= ------------------------------------------

p minusEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs -= rhs;
    assert lhs == expectedResult;
}

p minusEqualTestInnerUnsafe<TRhs>(int* lhs, const TRhs rhs, const int* expectedResult) {
    unsafe {
        lhs -= rhs;
    }
    assert lhs == expectedResult;
}

p minusEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    minusEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    minusEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    minusEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    minusEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p minusEqualTest() {
    // Lhs is double
    minusEqualTestOuter<double, double>(1.234, 98.7654, -97.5314, 97.5314, -99.9994, 99.9994);
    // Lhs is int
    minusEqualTestOuter<int, int>(78, 674, -596, 596, -752, 752);
    minusEqualTestOuter<int, short>(78, 7s, 71, -71, -85, 85);
    minusEqualTestOuter<int, long>(78, 2384723l, -2384645, 2384645, -2384801, 2384801);
    // Lhs is short
    minusEqualTestOuter<short, int>(78s, 674, -596s, 596s, -752s, 752s);
    minusEqualTestOuter<short, short>(78s, 7s, 71s, -71s, -85s, 85s);
    // Note: wrap-around consistent with short semantics
    minusEqualTestOuter<short, long>(78s, 2384723l, cast<short>(78s - 2384723l), cast<short>(-78s - -2384723l), cast<short>(-78s - 2384723l), cast<short>(78s - -2384723l));
    // Lhs is long
    minusEqualTestOuter<long, int>(78l, 674, -596l, 596l, -752l, 752l);
    minusEqualTestOuter<long, short>(78l, 7s, 71l, -71l, -85l, 85l);
    minusEqualTestOuter<long, long>(78l, 2384723l, -2384645l, 2384645l, -2384801l, 2384801l);
    // Lhs is char
    minusEqualTestInner<char, int>('A', 5, '<');
    minusEqualTestInner<char, int>('A', -5, 'F');
    // Lhs is ptr
    int[5] input = [0, 0, 0, 0, 0];
    minusEqualTestInnerUnsafe(&input[2], 2, &input[0]);
    minusEqualTestInnerUnsafe(&input[2], -2, &input[4]);
    minusEqualTestInnerUnsafe(&input[2], 2s, &input[0]);
    minusEqualTestInnerUnsafe(&input[2], -2s, &input[4]);
    minusEqualTestInnerUnsafe(&input[2], 2l, &input[0]);
    minusEqualTestInnerUnsafe(&input[2], -2l, &input[4]);
}

// ------------------------------------------ *= ------------------------------------------

p mulEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs *= rhs;
    assert lhs == expectedResult;
}

p mulEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    mulEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    mulEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    mulEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    mulEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p mulEqualTest() {
    // Lhs double
    mulEqualTestOuter<double, double>(1.5, 2.0, 3.0, 3.0, -3.0, -3.0);
    // Lhs int
    mulEqualTestOuter<int, int>(6, 7, 42, 42, -42, -42);
    mulEqualTestOuter<int, short>(6, 3s, 18, 18, -18, -18);
    mulEqualTestOuter<int, long>(6, 5l, 30, 30, -30, -30);
    // Lhs short
    mulEqualTestOuter<short, int>(6s, 7, 42s, 42s, -42s, -42s);
    mulEqualTestOuter<short, short>(6s, 3s, 18s, 18s, -18s, -18s);
    // Note: wrap-around consistent with short semantics
    mulEqualTestOuter<short, long>(200s, 2000l, cast<short>(200 * 2000), cast<short>(-200 * -2000), cast<short>(-200 * 2000), cast<short>(200 * -2000));
    // Lhs long
    mulEqualTestOuter<long, int>(6l, 7, 42l, 42l, -42l, -42l);
    mulEqualTestOuter<long, short>(6l, 3s, 18l, 18l, -18l, -18l);
    mulEqualTestOuter<long, long>(6l, 5l, 30l, 30l, -30l, -30l);
}

// ------------------------------------------ /= ------------------------------------------

p divEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs /= rhs;
    assert lhs == expectedResult;
}

p divEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    divEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    divEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    divEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    divEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p divEqualTest() {
    // Lhs double
    divEqualTestOuter<double, double>(9.0, 3.0, 3.0, 3.0, -3.0, -3.0);
    // Lhs int
    divEqualTestOuter<int, int>(42, 7, 6, 6, -6, -6);
    divEqualTestOuter<int, short>(42, 3s, 14, 14, -14, -14);
    divEqualTestOuter<int, long>(42, 6l, 7, 7, -7, -7);
    // Lhs short
    divEqualTestOuter<short, int>(42s, 7, 6s, 6s, -6s, -6s);
    divEqualTestOuter<short, short>(42s, 3s, 14s, 14s, -14s, -14s);
    divEqualTestOuter<short, long>(100s, 25l, 4s, 4s, -4s,- 4s);
    // Lhs long
    divEqualTestOuter<long, int>(42l, 7, 6l, 6l, -6l, -6l);
    divEqualTestOuter<long, short>(42l, 3s, 14l, 14l, -14l, -14l);
    divEqualTestOuter<long, long>(42l, 6l, 7l, 7l, -7l, -7l);
}

// ------------------------------------------ %= ------------------------------------------

p remEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs %= rhs;
    assert lhs == expectedResult;
}

p remEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2, const TLhs expectedResult3, const TLhs expectedResult4) {
    remEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    remEqualTestInner(-lhs, -rhs, expectedResult2); // Lhs -, Rhs -
    remEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    remEqualTestInner(lhs, -rhs, expectedResult4);  // Lhs +, Rhs -
}

p remEqualTest() {
    // Lhs double
    remEqualTestOuter<double, double>(9.0, 3.0, 0.0, 0.0, 0.0, 0.0);
    // Lhs int
    remEqualTestOuter<int, int>(42, 7, -0, -0, 0, 0);
    remEqualTestOuter<int, short>(42, 8s, 2, -2, -2, 2);
    remEqualTestOuter<int, long>(42, 9l, 6, -6, -6, 6);
    // Lhs short
    remEqualTestOuter<short, int>(42s, 7, -0s, -0s, 0s, 0s);
    remEqualTestOuter<short, short>(42s, 8s, 2s, -2s, -2s, 2s);
    remEqualTestOuter<short, long>(100s, 26l, 22s, -22s, -22s, 22s);
    // Lhs long
    remEqualTestOuter<long, int>(42l, 7, -0l, -0l, 0l, 0l);
    remEqualTestOuter<long, short>(42l, 10s, 2l, -2l, -2l, 2l);
    remEqualTestOuter<long, long>(10932847123l, 234324l, 226579l, -226579l, -226579l, 226579l);
    // Lhs byte
    remEqualTestInner<byte, byte>(cast<byte>(42), cast<byte>(41), cast<byte>(1));
}

// ------------------------------------------ <<= -----------------------------------------

p shlEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs <<= rhs;
    assert lhs == expectedResult;
}

p shlEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2) {
    shlEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    shlEqualTestInner(-lhs, rhs, expectedResult2);  // Lhs -, Rhs +
}

p shlEqualTest() {
    // Lhs int
    shlEqualTestOuter<int, int>(5, 3, 40, -40);
    shlEqualTestOuter<int, short>(5, 2s, 20, -20);
    shlEqualTestOuter<int, long>(5, 4l, 80, -80);
    // Lhs short
    shlEqualTestOuter<short, int>(8s, 2, 32s, -32s);
    shlEqualTestOuter<short, short>(8s, 1s, 16s, -16s);
    shlEqualTestOuter<short, long>(8s, 6l, 512s, -512s);
    // Lhs long
    shlEqualTestOuter<long, int>(7l, 7, 896l, -896l);
    shlEqualTestOuter<long, short>(7l, 10s, 7168l, -7168l);
    shlEqualTestOuter<long, long>(1234876l, 21l, 2589722673152l, -2589722673152l);
    // Lhs byte
    shlEqualTestInner<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(84));
}

// ------------------------------------------ >>= -----------------------------------------

p shrEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs >>= rhs;
    assert lhs == expectedResult;
}

p shrEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult1, const TLhs expectedResult2) {
    shrEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    shrEqualTestInner(-lhs, rhs, expectedResult2);  // Lhs -, Rhs +
}

p shrEqualTest() {
    // Lhs int
    shrEqualTestOuter<int, int>(5, 3, 0, -1);
    shrEqualTestOuter<int, short>(5, 2s, 1, -2);
    shrEqualTestOuter<int, long>(5, 1l, 2, -3);
    // Lhs short
    shrEqualTestOuter<short, int>(8s, 2, 2s, -2s);
    shrEqualTestOuter<short, short>(8s, 1s, 4s, 32764s);
    shrEqualTestOuter<short, long>(8s, 3l, 1s, -1s);
    // Lhs long
    shrEqualTestOuter<long, int>(23425l, 7, 183l, -184l);
    shrEqualTestOuter<long, short>(34587334534l, 10s, 33776693l, -33776694l);
    shrEqualTestOuter<long, long>(1234876l, 21l, 0l, -1l);
    // Lhs byte
    shrEqualTestInner<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(21));
}

// ------------------------------------------ &= ------------------------------------------

p andEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs &= rhs;
    assert lhs == expectedResult;
}

p andEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    andEqualTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p andEqualTest() {
    // Lhs int
    andEqualTestOuter<int, int>(5, 3, 1);
    andEqualTestOuter<int, short>(5, 2s, 0);
    andEqualTestOuter<int, long>(5, 1l, 1);
    // Lhs short
    andEqualTestOuter<short, int>(8s, 2, 0s);
    andEqualTestOuter<short, short>(8s, 1s, 0s);
    andEqualTestOuter<short, long>(8s, 3l, 0s);
    // Lhs long
    andEqualTestOuter<long, int>(23425l, 7, 1l);
    andEqualTestOuter<long, short>(34587334534l, 10s, 2l);
    andEqualTestOuter<long, long>(1234876l, 21l, 20l);
    // Lhs byte
    andEqualTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(0));
}

// ------------------------------------------ |= ------------------------------------------

p orEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs |= rhs;
    assert lhs == expectedResult;
}

p orEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    orEqualTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p orEqualTest() {
    // Lhs int
    orEqualTestOuter<int, int>(5, 3, 7);
    orEqualTestOuter<int, short>(5, 2s, 7);
    orEqualTestOuter<int, long>(5, 1l, 5);
    // Lhs short
    orEqualTestOuter<short, int>(8s, 2, 10s);
    orEqualTestOuter<short, short>(8s, 1s, 9s);
    orEqualTestOuter<short, long>(8s, 3l, 11s);
    // Lhs long
    orEqualTestOuter<long, int>(23425l, 7, 23431l);
    orEqualTestOuter<long, short>(34587334534l, 10s, 34587334542l);
    orEqualTestOuter<long, long>(1234876l, 21l, 1234877l);
    // Lhs byte
    orEqualTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(43));
}

// ------------------------------------------ ^= ------------------------------------------

p xorEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    lhs ^= rhs;
    assert lhs == expectedResult;
}

p xorEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    xorEqualTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p xorEqualTest() {
    // Lhs int
    xorEqualTestOuter<int, int>(5, 3, 6);
    xorEqualTestOuter<int, short>(5, 2s, 7);
    xorEqualTestOuter<int, long>(5, 1l, 4);
    // Lhs short
    xorEqualTestOuter<short, int>(8s, 2, 10s);
    xorEqualTestOuter<short, short>(8s, 1s, 9s);
    xorEqualTestOuter<short, long>(8s, 3l, 11s);
    // Lhs long
    xorEqualTestOuter<long, int>(23425l, 7, 23430l);
    xorEqualTestOuter<long, short>(34587334534l, 10s, 34587334540l);
    xorEqualTestOuter<long, long>(1234876l, 21l, 1234857l);
    // Lhs byte
    xorEqualTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(43));
}

// ------------------------------------------ ^ ------------------------------------------

p bitwiseXorTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs ^ rhs;
    assert actualResult == expectedResult;
}

p bitwiseXorTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    bitwiseXorTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p bitwiseXorTest() {
    // Lhs int
    bitwiseXorTestOuter<int, int>(5, 3, 6);
    // Lhs short
    bitwiseXorTestOuter<short, short>(8s, 1s, 9s);
    // Lhs long
    bitwiseXorTestOuter<long, long>(1234876l, 21l, 1234857l);
    // Lhs byte
    bitwiseXorTestOuter<byte, byte>(cast<byte>(15), cast<byte>(23), cast<byte>(24));
    // Lhs bool
    bitwiseXorTestOuter<bool, bool>(false, false, false);
    bitwiseXorTestOuter<bool, bool>(false, true, true);
    bitwiseXorTestOuter<bool, bool>(true, false, true);
    bitwiseXorTestOuter<bool, bool>(true, true, false);
}

// ------------------------------------------ | ------------------------------------------

p bitwiseOrTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs | rhs;
    assert actualResult == expectedResult;
}

p bitwiseOrTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    bitwiseOrTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p bitwiseOrTest() {
    // Lhs int
    bitwiseOrTestOuter<int, int>(5, 3, 7);
    // Lhs short
    bitwiseOrTestOuter<short, short>(8s, 1s, 9s);
    // Lhs long
    bitwiseOrTestOuter<long, long>(1234876l, 21l, 1234877l);
    // Lhs byte
    bitwiseOrTestOuter<byte, byte>(cast<byte>(42), cast<byte>(1), cast<byte>(43));
    // Lhs bool
    bitwiseOrTestOuter<bool, bool>(false, false, false);
    bitwiseOrTestOuter<bool, bool>(false, true, true);
    bitwiseOrTestOuter<bool, bool>(true, false, true);
    bitwiseOrTestOuter<bool, bool>(true, true, true);
}

// ------------------------------------------ & ------------------------------------------

p bitwiseAndTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    const TLhs actualResult = lhs & rhs;
    assert actualResult == expectedResult;
}

p bitwiseAndTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const TLhs expectedResult) {
    bitwiseAndTestInner(lhs, rhs, expectedResult);   // Lhs +, Rhs +
}

p bitwiseAndTest() {
    // Lhs int
    bitwiseAndTestOuter<int, int>(5, 3, 1);
    // Lhs short
    bitwiseAndTestOuter<short, short>(8s, 1s, 0s);
    // Lhs long
    bitwiseAndTestOuter<long, long>(1234876l, 21l, 20l);
    // Lhs byte
    bitwiseAndTestOuter<byte, byte>(cast<byte>(15), cast<byte>(23), cast<byte>(7));
    // Lhs bool
    bitwiseAndTestOuter<bool, bool>(false, false, false);
    bitwiseAndTestOuter<bool, bool>(false, true, false);
    bitwiseAndTestOuter<bool, bool>(true, false, false);
    bitwiseAndTestOuter<bool, bool>(true, true, true);
}

// ------------------------------------------ == -----------------------------------------

p equalTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs == rhs;
    assert actualResult == expectedResult;
}

p equalTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    equalTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    equalTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    equalTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    equalTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p equalTest() {
    // Lhs is ptr
    int i = 213;
    int* iPtr = &i;
    equalTestInner<int*, int*>(iPtr, iPtr, false);
    // Lhs double
    equalTestOuter<double, int>(87.0, 87, true, false, false, true);
    equalTestOuter<double, short>(14.0, 14s, true, false, false, true);
    equalTestOuter<double, long>(2349234.0, 2349234l, true, false, false, true);
    // Lhs int
    equalTestOuter<int, double>(12345, 12345.0, true, false, false, true);
    equalTestOuter<int, int>(5, 5, true, false, false, true);
    equalTestOuter<int, short>(-234, -234s, true, false, false, true);
    equalTestOuter<int, long>(-9999999, 9999999l, false, true, true, false);
    equalTestInner<int, char>(67, 'C', true);
    // Lhs short
    equalTestOuter<short, double>(12345s, 12345.0, true, false, false, true);
    equalTestOuter<short, int>(5s, 5, true, false, false, true);
    equalTestOuter<short, short>(-234s, -234s, true, false, false, true);
    equalTestOuter<short, long>(-999s, 999l, false, true, true, false);
    equalTestInner<short, char>(68s, 'D', true);
    // Lhs long
    equalTestOuter<long, double>(12345l, 12345.0, true, false, false, true);
    equalTestOuter<long, int>(5l, 5, true, false, false, true);
    equalTestOuter<long, short>(-234l, -234s, true, false, false, true);
    equalTestOuter<long, long>(-999l, 999l, false, true, true, false);
    equalTestInner<long, char>(68l, 'D', true);
    // Lhs byte
    equalTestInner<byte, byte>(cast<byte>(15), cast<byte>(15), true);
    // Lhs char
    equalTestInner<char, int>('x', -15, false);
    equalTestInner<char, short>('5', 53s, true);
    equalTestInner<char, long>('+', 43l, true);
    equalTestInner<char, char>('#', '#', true);
    // Lhs string
    equalTestInner<string, string>("this is a test", "this is a test", true);
    equalTestInner<string, string>("string", "strong", false);
    String strA = String("this is a test");
    String strB = String("strong");
    equalTestInner<string, string>("this is a test", strA.getRaw(), true);
    equalTestInner<string, string>("string", strB.getRaw(), false);
    // Lhs bool
    equalTestInner<bool, bool>(false, false, false);
    equalTestInner<bool, bool>(false, true, true);
    equalTestInner<bool, bool>(true, false, true);
    equalTestInner<bool, bool>(true, true, false);
    // Lhs function
    const dyn funcA = f<int>(bool b, double d) { return 123; };
    const dyn funcB = f<int>(bool b, double d) { return 456; };
    equalTestInner<f<int>(bool, double), f<int>(bool, double)>(funcA, funcA, true);
    equalTestInner<f<int>(bool, double), f<int>(bool, double)>(funcA, funcB, false);
    // Lhs procedure
    const dyn procA = p(string s, char c) {};
    const dyn procB = p(string s, char c) {};
    equalTestInner<p(string, char), p(string, char)>(procA, procA, true);
    equalTestInner<p(string, char), p(string, char)>(procA, procB, false);
}

// ------------------------------------------ != -----------------------------------------

p notEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs == rhs;
    assert actualResult == expectedResult;
}

p notEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    notEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    notEqualTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    notEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    notEqualTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p notEqualTest() {
    // Lhs is ptr
    int i = 213;
    int* iPtr = &i;
    notEqualTestInner<int*, int*>(iPtr, iPtr, true);
    // Lhs double
    notEqualTestOuter<double, int>(87.0, 87, false, true, true, false);
    notEqualTestOuter<double, short>(14.0, 14s, false, true, true, false);
    notEqualTestOuter<double, long>(2349234.0, 2349234l, false, true, true, false);
    // Lhs int
    notEqualTestOuter<int, double>(12345, 12345.0, false, true, true, false);
    notEqualTestOuter<int, int>(5, 5, false, true, true, false);
    notEqualTestOuter<int, short>(-234, -234s, false, true, true, false);
    notEqualTestOuter<int, long>(-9999999, 9999999l, true, false, false, true);
    notEqualTestInner<int, char>(67, 'C', false);
    // Lhs short
    notEqualTestOuter<short, double>(12345s, 12345.0, false, true, true, false);
    notEqualTestOuter<short, int>(5s, 5, false, true, true, false);
    notEqualTestOuter<short, short>(-234s, -234s, false, true, true, false);
    notEqualTestOuter<short, long>(-999s, 999l, true, false, false, true);
    notEqualTestInner<short, char>(68s, 'D', false);
    // Lhs long
    notEqualTestOuter<long, double>(12345l, 12345.0, false, true, true, false);
    notEqualTestOuter<long, int>(5l, 5, false, true, true, false);
    notEqualTestOuter<long, short>(-234l, -234s, false, true, true, false);
    notEqualTestOuter<long, long>(-999l, 999l, true, false, false, true);
    notEqualTestInner<long, char>(68l, 'D', false);
    // Lhs byte
    notEqualTestInner<byte, byte>(cast<byte>(15), cast<byte>(15), false);
    // Lhs char
    notEqualTestInner<char, int>('x', -15, true);
    notEqualTestInner<char, short>('5', 53s, false);
    notEqualTestInner<char, long>('+', 43l, false);
    notEqualTestInner<char, char>('#', '#', false);
    // Lhs string
    notEqualTestInner<string, string>("this is a test", "this is a test", false);
    notEqualTestInner<string, string>("string", "strong", true);
    String strA = String("this is a test");
    String strB = String("strong");
    notEqualTestInner<string, string>("this is a test", strA.getRaw(), false);
    notEqualTestInner<string, string>("string", strB.getRaw(), true);
    // Lhs bool
    notEqualTestInner<bool, bool>(false, false, true);
    notEqualTestInner<bool, bool>(false, true, false);
    notEqualTestInner<bool, bool>(true, false, false);
    notEqualTestInner<bool, bool>(true, true, true);
    // Lhs function
    const dyn funcA = f<int>(bool b, double d) { return 123; };
    const dyn funcB = f<int>(bool b, double d) { return 456; };
    notEqualTestInner<f<int>(bool, double), f<int>(bool, double)>(funcA, funcA, false);
    notEqualTestInner<f<int>(bool, double), f<int>(bool, double)>(funcA, funcB, true);
    // Lhs procedure
    const dyn procA = p(string s, char c) {};
    const dyn procB = p(string s, char c) {};
    notEqualTestInner<p(string, char), p(string, char)>(procA, procA, false);
    notEqualTestInner<p(string, char), p(string, char)>(procA, procB, true);
}

// ------------------------------------------ < ------------------------------------------

p lessTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs < rhs;
    assert actualResult == expectedResult;
}

p lessTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    lessTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    lessTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    lessTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    lessTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p lessTest() {
    // Lhs double
    lessTestOuter<double, double>(87.123, 87.124, true, false, false, true);
    lessTestOuter<double, int>(87.0, 88, true, false, false, true);
    lessTestOuter<double, short>(14.0, 15s, true, false, false, true);
    lessTestOuter<double, long>(2349234.0, 2349235l, true, false, false, true);
    // Lhs int
    lessTestOuter<int, double>(12345, 12345.1, true, false, false, true);
    lessTestOuter<int, int>(5, 6, true, false, false, true);
    lessTestOuter<int, short>(-234, -233s, true, false, false, true);
    lessTestOuter<int, long>(9999999, -9999999l, false, true, true, false);
    // Lhs short
    lessTestOuter<short, double>(12345s, 12345.423, true, false, false, true);
    lessTestOuter<short, int>(5s, 6, true, false, false, true);
    lessTestOuter<short, short>(-234s, -233s, true, false, false, true);
    lessTestOuter<short, long>(999s, -999l, false, true, true, false);
    // Lhs long
    lessTestOuter<long, double>(12345l, 12345.1, true, false, false, true);
    lessTestOuter<long, int>(5l, 6, true, false, false, true);
    lessTestOuter<long, short>(-234l, -233s, true, false, false, true);
    lessTestOuter<long, long>(999l, -999l, false, true, true, false);
    // Lhs byte
    lessTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), true);
    // Lhs char
    lessTestInner<char, char>('#', '#', false);
}

// ------------------------------------------ > ------------------------------------------

p greaterTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs > rhs;
    assert actualResult == expectedResult;
}

p greaterTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    greaterTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    greaterTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    greaterTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    greaterTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p greaterTest() {
    // Lhs double
    greaterTestOuter<double, double>(87.123, 87.124, false, true, true, false);
    greaterTestOuter<double, int>(87.0, 88, false, true, true, false);
    greaterTestOuter<double, short>(14.0, 15s, false, true, true, false);
    greaterTestOuter<double, long>(2349234.0, 2349235l, false, true, true, false);
    // Lhs int
    greaterTestOuter<int, double>(12345, 12345.1, false, true, true, false);
    greaterTestOuter<int, int>(5, 6, false, true, true, false);
    greaterTestOuter<int, short>(-234, -233s, false, true, true, false);
    greaterTestOuter<int, long>(9999999, -9999999l, true, false, false, true);
    // Lhs short
    greaterTestOuter<short, double>(12345s, 12345.423, false, true, true, false);
    greaterTestOuter<short, int>(5s, 6, false, true, true, false);
    greaterTestOuter<short, short>(-234s, -233s, false, true, true, false);
    greaterTestOuter<short, long>(999s, -999l, true, false, false, true);
    // Lhs long
    greaterTestOuter<long, double>(12345l, 12345.1, false, true, true, false);
    greaterTestOuter<long, int>(5l, 6, false, true, true, false);
    greaterTestOuter<long, short>(-234l, -233s, false, true, true, false);
    greaterTestOuter<long, long>(999l, -999l, true, false, false, true);
    // Lhs byte
    greaterTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), false);
    // Lhs char
    greaterTestInner<char, char>('#', '#', false);
}

// ------------------------------------------ <= -----------------------------------------

p lessEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs <= rhs;
    assert actualResult == expectedResult;
}

p lessEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    lessEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    lessEqualTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    lessEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    lessEqualTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p lessEqualTest() {
    // Lhs double
    lessEqualTestOuter<double, double>(87.123, 87.124, true, false, false, true);
    lessEqualTestOuter<double, int>(87.0, 88, true, false, false, true);
    lessEqualTestOuter<double, short>(14.0, 15s, true, false, false, true);
    lessEqualTestOuter<double, long>(2349234.0, 2349235l, true, false, false, true);
    // Lhs int
    lessEqualTestOuter<int, double>(12345, 12345.1, true, false, false, true);
    lessEqualTestOuter<int, int>(5, 6, true, false, false, true);
    lessEqualTestOuter<int, short>(-234, -233s, true, false, false, true);
    lessEqualTestOuter<int, long>(9999999, -9999999l, false, true, true, false);
    // Lhs short
    lessEqualTestOuter<short, double>(12345s, 12345.423, true, false, false, true);
    lessEqualTestOuter<short, int>(5s, 6, true, false, false, true);
    lessEqualTestOuter<short, short>(-234s, -233s, true, false, false, true);
    lessEqualTestOuter<short, long>(999s, -999l, false, true, true, false);
    // Lhs long
    lessEqualTestOuter<long, double>(12345l, 12345.1, true, false, false, true);
    lessEqualTestOuter<long, int>(5l, 6, true, false, false, true);
    lessEqualTestOuter<long, short>(-234l, -233s, true, false, false, true);
    lessEqualTestOuter<long, long>(999l, -999l, false, true, true, false);
    // Lhs byte
    lessEqualTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), true);
    // Lhs char
    lessEqualTestInner<char, char>('#', '#', true);
}

// ------------------------------------------ >= -----------------------------------------

p greaterEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs >= rhs;
    assert actualResult == expectedResult;
}

p greaterEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    greaterEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    greaterEqualTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    greaterEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    greaterEqualTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p greaterEqualTest() {
    // Lhs double
    greaterEqualTestOuter<double, double>(87.123, 87.124, false, true, true, false);
    greaterEqualTestOuter<double, int>(87.0, 88, false, true, true, false);
    greaterEqualTestOuter<double, short>(14.0, 15s, false, true, true, false);
    greaterEqualTestOuter<double, long>(2349234.0, 2349235l, false, true, true, false);
    // Lhs int
    greaterEqualTestOuter<int, double>(12345, 12345.1, false, true, true, false);
    greaterEqualTestOuter<int, int>(5, 6, false, true, true, false);
    greaterEqualTestOuter<int, short>(-234, -233s, false, true, true, false);
    greaterEqualTestOuter<int, long>(9999999, -9999999l, true, false, false, true);
    // Lhs short
    greaterEqualTestOuter<short, double>(12345s, 12345.423, false, true, true, false);
    greaterEqualTestOuter<short, int>(5s, 6, false, true, true, false);
    greaterEqualTestOuter<short, short>(-234s, -233s, false, true, true, false);
    greaterEqualTestOuter<short, long>(999s, -999l, true, false, false, true);
    // Lhs long
    greaterEqualTestOuter<long, double>(12345l, 12345.1, false, true, true, false);
    greaterEqualTestOuter<long, int>(5l, 6, false, true, true, false);
    greaterEqualTestOuter<long, short>(-234l, -233s, false, true, true, false);
    greaterEqualTestOuter<long, long>(999l, -999l, true, false, false, true);
    // Lhs byte
    greaterEqualTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), false);
    // Lhs char
    greaterEqualTestInner<char, char>('#', '#', true);
}

f<int> main() {
    plusEqualTest();    // +=
    minusEqualTest();   // -=
    mulEqualTest();     // *=
    divEqualTest();     // /=
    remEqualTest();     // %=
    shlEqualTest();     // <<=
    shrEqualTest();     // >>=
    andEqualTest();     // &=
    orEqualTest();      // |=
    xorEqualTest();     // ^=
    bitwiseOrTest();    // |
    bitwiseXorTest();   // ^
    bitwiseAndTest();   // &
    equalTest();        // ==
    notEqualTest();     // !=
    lessTest();         // <
    greaterTest();      // >
    lessEqualTest();    // >
    greaterEqualTest(); // >
    // ToDo: Extend

    printf("All assertions passed!");
}