import "std/io/file";

f<int> main() {
    // Write file
    Result<File> fileResult = openFile("./test-file.txt", MODE_WRITE);
    assert fileResult.isOk();
    File file = fileResult.unwrap();
    bool _ = file.write("Hello, world!\n");
    _ = file.close();

    // Read file
    fileResult = openFile("./test-file.txt", MODE_READ);
    assert fileResult.isOk();
    file = fileResult.unwrap();
    assert file.readLine() == String("Hello, world!");
    _ = file.close();

    // Append file
    fileResult = openFile("./test-file.txt", MODE_APPEND);
    assert fileResult.isOk();
    file = fileResult.unwrap();
    _ = file.write("Hello, again!\n");
    _ = file.close();

    // Read file
    fileResult = openFile("./test-file.txt", MODE_READ);
    assert fileResult.isOk();
    file = fileResult.unwrap();
    assert file.readLine() == String("Hello, world!");
    assert file.readLine() == String("Hello, again!");
    _ = file.close();

    printf("All assertions passed!");
}