import "std/test/lifetime-object";

f<LifetimeObject> spawnLO() {
    return LifetimeObject();
}

f<LifetimeObject> decideOnLOConstRef(bool cond, const LifetimeObject& lo1, const LifetimeObject& lo2) {
    cond ? lo1 : lo2; // Should not do a copy
    LifetimeObject loCopy = cond ? lo1 : lo2; // Shoud do a copy
    const LifetimeObject& loRef = cond ? lo1 : lo2; // Should not do a copy
    return cond ? lo1 : lo2; // Return statement should do a copy
}

f<LifetimeObject> decideOnLORef(bool cond, LifetimeObject& lo1, LifetimeObject& lo2) {
    cond ? lo1 : lo2; // Should not do a copy
    LifetimeObject loCopy = cond ? lo1 : lo2; // Shoud do a copy
    const LifetimeObject& loRef = cond ? lo1 : lo2; // Should not do a copy
    return cond ? lo1 : lo2; // Return statement should do a copy
}

f<LifetimeObject> decideOnLOVal(bool cond, LifetimeObject lo1, LifetimeObject lo2) {
    cond ? lo1 : lo2; // Shoud do a copy, although the result is ignored
    LifetimeObject loCopy = cond ? lo1 : lo2; // Shoud do a copy
    const LifetimeObject& loRef = cond ? lo1 : lo2; // Should do a copy
    return cond ? lo1 : lo2; // Return statement should do a copy
}

f<int> main() {
    // Ignored return value of ctor
    printf("Ignored return value of ctor:\n");
    {
        LifetimeObject();
    }

    // Normal lifecycle
    printf("Normal lifecycle:\n");
    {
        LifetimeObject lo = LifetimeObject(); // ctor call
        LifetimeObject loCopy = lo; // copy ctor call
    }

    // Return from lambda as value
    printf("Return from lambda as value:\n");
    {
        const f<LifetimeObject>() spawnLO = f<LifetimeObject>() {
            return LifetimeObject();
        };

        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    // Return from lambda as reference
    printf("Return from lambda as reference:\n");
    {
        LifetimeObject loOrig = LifetimeObject();
        const f<LifetimeObject&>() spawnLO = f<LifetimeObject&>() {
            return loOrig;
        };

        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Copy
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    // Return from lambda as const reference
    printf("Return from lambda as const reference:\n");
    {
        LifetimeObject loOrig = LifetimeObject();
        const f<const LifetimeObject&>() spawnLO = f<const LifetimeObject&>() {
            return loOrig;
        };

        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Copy
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    // Return from function as value
    printf("Return from function as value:\n");
    {
        // No return value receiver
        spawnLO(); // Anonymous symbol
        // Return value receiver - value
        LifetimeObject lo = spawnLO(); // Assigned to lo
        // Return value receiver - const ref
        const LifetimeObject& loConstRef = spawnLO(); // Assigned to loConstRef
    }

    printf("Ternary (true temporary, false temporary)\n");
    {
        bool cond = true;
        LifetimeObject loCopy1 = cond ? LifetimeObject() : LifetimeObject(); // ctor calls in both branches
        LifetimeObject loCopy2 = !cond ? LifetimeObject() : LifetimeObject(); // ctor calls in both branches
    }

    printf("Ternary (true temporary, false not temporary)\n");
    {
        bool cond = true;
        LifetimeObject lo = LifetimeObject();
        LifetimeObject loCopy1 = cond ? LifetimeObject() : lo; // ctor in true branch, copy ctor in false branch
        LifetimeObject loCopy2 = !cond ? LifetimeObject() : lo; // ctor in true branch, copy ctor in false branch
    }

    printf("Ternary (true not temporary, false temporary)\n");
    {
        bool cond = true;
        LifetimeObject lo = LifetimeObject();
        LifetimeObject loCopy1 = cond ? lo : LifetimeObject(); // copy ctor in true branch, ctor in false branch
        LifetimeObject loCopy2 = !cond ? lo : LifetimeObject(); // copy ctor in true branch, ctor in false branch
    }

    printf("Ternary (true not temporary, false not temporary)\n");
    {
        bool cond = true;
        LifetimeObject lo1 = LifetimeObject();
        LifetimeObject lo2 = LifetimeObject();
        LifetimeObject loCopy1 = cond ? lo1 : lo2; // copy ctor call in both branches
        LifetimeObject loCopy2 = !cond ? lo1 : lo2; // copy ctor call in both branches
    }

    printf("Ternary function (const ref) return:\n");
    {
        bool cond = true;
        LifetimeObject lo1 = LifetimeObject();
        LifetimeObject lo2 = LifetimeObject();
        LifetimeObject lo3 = decideOnLOConstRef(cond, lo1, lo2);
        LifetimeObject lo4 = decideOnLOConstRef(!cond, lo1, lo2);
    }

    printf("Ternary function (ref) return:\n");
    {
        bool cond = true;
        LifetimeObject lo1 = LifetimeObject();
        LifetimeObject lo2 = LifetimeObject();
        LifetimeObject lo3 = decideOnLORef(cond, lo1, lo2);
        LifetimeObject lo4 = decideOnLORef(!cond, lo1, lo2);
    }

    printf("Ternary function (val) return:\n");
    {
        bool cond = true;
        LifetimeObject lo1 = LifetimeObject();
        LifetimeObject lo2 = LifetimeObject();
        LifetimeObject lo3 = decideOnLOVal(cond, lo1, lo2);
        LifetimeObject lo4 = decideOnLOVal(!cond, lo1, lo2);
    }

    printf("Ternary receiving function result:\n");
    {
        bool cond = false;
        LifetimeObject lo1 = cond ? spawnLO() : spawnLO();
        LifetimeObject lo2 = !cond ? (cond ? spawnLO() : spawnLO()) : spawnLO();
    }
}