// TEST: --sanitizer=address -g

f<int> main() {
    heap int* iPtr = sNew<int>();
    *iPtr = 123;
    unsafe {
        sDealloc(cast<heap byte*>(iPtr));
    }
    *iPtr = 321;
}