type TLhs dyn;
type TRhs dyn;

// ------------------------------------------ <= -----------------------------------------

p lessEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs <= rhs;
    assert actualResult == expectedResult;
}

p lessEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    lessEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    lessEqualTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    lessEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    lessEqualTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p lessEqualTest() {
    // Lhs double
    lessEqualTestOuter<double, double>(87.123, 87.124, true, false, false, true);
    lessEqualTestOuter<double, int>(87.0, 88, true, false, false, true);
    lessEqualTestOuter<double, short>(14.0, 15s, true, false, false, true);
    lessEqualTestOuter<double, long>(2349234.0, 2349235l, true, false, false, true);
    // Lhs int
    lessEqualTestOuter<int, double>(12345, 12345.1, true, false, false, true);
    lessEqualTestOuter<int, int>(5, 6, true, false, false, true);
    lessEqualTestOuter<int, short>(-234, -233s, true, false, false, true);
    lessEqualTestOuter<int, long>(9999999, -9999999l, false, true, true, false);
    // Lhs short
    lessEqualTestOuter<short, double>(12345s, 12345.423, true, false, false, true);
    lessEqualTestOuter<short, int>(5s, 6, true, false, false, true);
    lessEqualTestOuter<short, short>(-234s, -233s, true, false, false, true);
    lessEqualTestOuter<short, long>(999s, -999l, false, true, true, false);
    // Lhs long
    lessEqualTestOuter<long, double>(12345l, 12345.1, true, false, false, true);
    lessEqualTestOuter<long, int>(5l, 6, true, false, false, true);
    lessEqualTestOuter<long, short>(-234l, -233s, true, false, false, true);
    lessEqualTestOuter<long, long>(999l, -999l, false, true, true, false);
    // Lhs byte
    lessEqualTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), true);
    // Lhs char
    lessEqualTestInner<char, char>('#', '#', true);
}

// ------------------------------------------ >= -----------------------------------------

p greaterEqualTestInner<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult) {
    const bool actualResult = lhs >= rhs;
    assert actualResult == expectedResult;
}

p greaterEqualTestOuter<TLhs, TRhs>(TLhs lhs, const TRhs rhs, const bool expectedResult1, const bool expectedResult2, const bool expectedResult3, const bool expectedResult4) {
    greaterEqualTestInner(lhs, rhs, expectedResult1);   // Lhs +, Rhs +
    greaterEqualTestInner(lhs, -rhs, expectedResult2);  // Lhs +, Rhs -
    greaterEqualTestInner(-lhs, rhs, expectedResult3);  // Lhs -, Rhs +
    greaterEqualTestInner(-lhs, -rhs, expectedResult4); // Lhs -, Rhs -
}

p greaterEqualTest() {
    // Lhs double
    greaterEqualTestOuter<double, double>(87.123, 87.124, false, true, true, false);
    greaterEqualTestOuter<double, int>(87.0, 88, false, true, true, false);
    greaterEqualTestOuter<double, short>(14.0, 15s, false, true, true, false);
    greaterEqualTestOuter<double, long>(2349234.0, 2349235l, false, true, true, false);
    // Lhs int
    greaterEqualTestOuter<int, double>(12345, 12345.1, false, true, true, false);
    greaterEqualTestOuter<int, int>(5, 6, false, true, true, false);
    greaterEqualTestOuter<int, short>(-234, -233s, false, true, true, false);
    greaterEqualTestOuter<int, long>(9999999, -9999999l, true, false, false, true);
    // Lhs short
    greaterEqualTestOuter<short, double>(12345s, 12345.423, false, true, true, false);
    greaterEqualTestOuter<short, int>(5s, 6, false, true, true, false);
    greaterEqualTestOuter<short, short>(-234s, -233s, false, true, true, false);
    greaterEqualTestOuter<short, long>(999s, -999l, true, false, false, true);
    // Lhs long
    greaterEqualTestOuter<long, double>(12345l, 12345.1, false, true, true, false);
    greaterEqualTestOuter<long, int>(5l, 6, false, true, true, false);
    greaterEqualTestOuter<long, short>(-234l, -233s, false, true, true, false);
    greaterEqualTestOuter<long, long>(999l, -999l, true, false, false, true);
    // Lhs byte
    greaterEqualTestInner<byte, byte>(cast<byte>(15), cast<byte>(16), false);
    // Lhs char
    greaterEqualTestInner<char, char>('#', '#', true);
}

f<int> main() {
    lessEqualTest(); // <=
    greaterEqualTest(); // >=
    // ToDo: Extend

    printf("All assertions passed!");
}