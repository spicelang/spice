type TestStruct struct {
    bool _f1
    int& f2
}

f<int> main() {
    int t = 123;
    dyn ts = TestStruct { true, t };
    printf("Before: %d\n", ts.f2);
    ts.f2++;
    printf("After: %d", t);
}