type T int;

f<int> main() {}