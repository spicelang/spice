/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/data/vector" as vector;

f<int> main() {
    dyn v = vector.Vector<int>{};
    v.push(4);
    v.push(2);
}*/

type T dyn;

public type Vector<T> struct {
    T* contents
    unsigned long capacity
    unsigned long size
    unsigned int itemSize
}

public f<int> Vector.get(long index) {
    if (index <= size) { // Note 'size' instead 'this.size'
        return 1;
    }
    return 0;
}

f<int> main() {
    dyn v = Vector<int>{};
    int v0 = v.get(0l);
}