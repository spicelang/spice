f<int> main() {
    /*if (true) {
        return 1;
    }
    while (true) {
        return 2;
    }*/
    printf("Test");
    return 0;
}