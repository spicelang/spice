import "os-test3";