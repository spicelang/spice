const int GLOBAL_TEST_VAR = 123;