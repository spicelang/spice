ext f<int> exteralFunction(dyn, int);

f<int> main() {
    extFunction(1, 3);
}