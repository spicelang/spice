type Test struct {
    int t
}

p Test.dtor() {
    printf("Dtor called!");
}

f<Test> test() {
    return Test{123};
}

f<int> main() {
   Test t = test();
   printf("%d", t.t);
}