/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*p testProc(int[]** nums) {
    int[] nums1 = **nums;
    //printf("De-referenced: %p\n", nums1);
    nums1[2] = 10;
    printf("1: %d\n", nums1[0]);
    printf("2: %d\n", nums1[1]);
    printf("3: %d\n", nums1[2]);
    printf("4: %d\n", nums1[3]);
}*/

f<int> main() {
    //int[4] intArray = { 1, 2, 3, 4 };
    //printf("1: %d\n", intArray[2]);
    //printf("Pointer: %p\n", intArray);
    //testProc(&&intArray);

    string test = "test";
    char c1 = test[2];
    printf("Char: %c\n", c1);
}