import "std/data/map";

f<int> main() {
    Map<int, string> map;
    assert map.getSize() == 0l;
    assert map.isEmpty();
    map.insert(1, "Hello");
    assert map.getSize() == 1l;
    assert !map.isEmpty();
    map.insert(2, "World");
    assert map.getSize() == 2l;
    map.insert(3, "Foo");
    assert map.getSize() == 3l;
    map.insert(4, "Bar");
    assert map.getSize() == 4l;
    assert map.contains(1);
    assert map.contains(2);
    assert map.contains(3);
    assert map.contains(4);
    assert map.get(1) == "Hello";
    assert map.get(2) == "World";
    assert map.get(3) == "Foo";
    assert map.get(4) == "Bar";
    map.remove(2);
    assert map.getSize() == 3l;
    assert !map.contains(2);
    assert !map.isEmpty();
    map.remove(1);
    assert map.getSize() == 2l;
    assert !map.contains(1);
    assert !map.isEmpty();
    string& foo = map.get(3);
    assert foo == "Foo";
    foo = "Baz";
    assert map.get(3) == "Baz";
    Result<string> bar = map.getSafe(4);
    assert bar.isOk();
    assert bar.unwrap() == "Bar";
    Result<string> baz = map.getSafe(5);
    assert baz.isErr();
    map.remove(3);
    assert map.getSize() == 1l;
    assert !map.contains(3);
    assert !map.isEmpty();
    map.remove(4);
    assert map.getSize() == 0l;
    assert !map.contains(4);
    assert map.isEmpty();
    printf("All assertions passed!\n");
}

/*import "std/os/env";
import "std/io/filepath";
import "bootstrap/ast/ast-nodes";
import "bootstrap/lexer/lexer";
import "bootstrap/parser/parser";

f<int> main() {
    String filePathString = getEnv("SPICE_STD_DIR") + "/../test/test-files/bootstrap-compiler/standalone-parser-test/test-file.spice";
    FilePath filePath = FilePath(filePathString);
    Lexer lexer = Lexer(filePath);
    Parser parser = Parser(lexer);
    ASTEntryNode* ast = parser.parse();
    assert ast != nil<ASTEntryNode*>;
    printf("All assertions passed!\n");
}*/