f<int> main() {
    string food = "Pizza";
    string* ptr = &food;

    printf("Pointer address: %p, value: %s", ptr, *ptr);

    dyn restoredFood = *ptr;
    printf("Restored value: %s", restoredFood);

    printf("Restored value address: %p", &restoredFood);
}