f<int> main() {
    int value = 1;
    value <<= 30;
    printf("Shifted value: %d", value);
}