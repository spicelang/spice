f<int> main() {
    while 5.6 {
        printf("Test");
    }
    return 0;
}