f<int> main() {
    string test = "Hello World!";
    string* testPtr = &test;
    *testPtr = "Hello Spice users!";
    printf("Value1: %s, pointer: %p, value: %s", test, testPtr, *testPtr);
}