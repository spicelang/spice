import "std/data/triple" as triple;

f<int> main() {
    triple::Triple<string, int, bool> stringIntBoolTriple = triple::Triple<string, int, bool>("Test", 1234, true);
    printf("First: %s\n", stringIntBoolTriple.getFirst());
    printf("Second: %d\n", stringIntBoolTriple.getSecond());
    printf("Third: %d\n", stringIntBoolTriple.getThird());
}