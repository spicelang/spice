//import "std/iterator/number-iterator";
import "std/runtime/iterator_rt";

f<int> main() {
    /*foreach int i : range(1, 5) {
        printf("%d\n", i);
    }*/

    Vector<int> vi = Vector<int>();
    vi.pushBack(123);
    vi.pushBack(4321);
    printf("Item 1: %d\n", vi.get(0));
    printf("Item 2: %d\n", vi.get(1));
    dyn it = iterate(vi);
    //printf("Get: %d\n", it.get());
    /*foreach int i : it {
        printf("Item: %d\n", i);
    }*/
}