/*import "std/data/queue" as que;

f<int> main() {
    dyn q1 = que.Queue<char>();
    q1.push('H');
    q1.push('e');
    q1.push('l');
    q1.push('l');
    q1.push('o');
    q1.push('!');
    printf("Size: %d, Capacity: %d\n", q1.getSize(), q1.getCapacity());
    while (!q1.isEmpty()) {
        printf("%c", q1.pop());
    }
    q1.dtor();
}*/

type T int|double|short|long;
type U bool[]|int[];

f<int> sumNumbers<T>(T[] numberArray, int arrayLength) {
    result = 0;
    for int i = 0; i < arrayLength; i++ {
        result += numberArray[i];
    }
}

p printData<U>(int arrayLength, U list) {
    for int i = 0; i < arrayLength; i++ {
        printf("Data: %d\n", list[i]);
    }
}

f<int> main() {
    short[7] numberList1 = { 1s, 2s, 3s, 4s, 5s, 6s, 7s };
    int result1 = sumNumbers(numberList1, len(numberList1));

    long[4] numberList2 = { 10l, 12l, 14l, 16l };
    int result2 = sumNumbers(numberList2, len(numberList2));

    dyn resultList = {result1, result2};
    printData(len(resultList), resultList);

    printf("Results: %d, %d\n", result1, result2);
}