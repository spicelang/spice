public type Test struct {
    public int u
}