f<int> main() {
    String test = String("Dies ist ein Test");
    char c = test[13l];
    printf("%s, %c", test, c);
}