type Test struct {
    int f1
    int f2
}

f<int> main() {
    int t = 123;
    switch (t) {
        case 1: {
            printf("1");
        }
        case Test: {
            printf("t");
        }
    }
}

/*import "std/data/optional";
import "std/data/stack";

f<int> main() {
    Stack<double> doubleStack = Stack<double>();
    doubleStack.push(4.566);

    dyn oi = Optional<Stack<double>>();
    printf("%d\n", oi.isPresent());
    oi.set(doubleStack);
    printf("%d\n", oi.isPresent());
    dyn res = oi.get();
    printf("%d\n", res.getSize());
    oi.clear();
    printf("%d\n", oi.isPresent());

    dyn oi2 = Optional<String>(String("This is a test"));
    assert oi2.isPresent();
}*/