import "std/iterators/number-iterator";
//import "std/iterators/array-iterator";

// Generic type definitions
type Numeric int|long|short;
type I dyn;

/**
 * Convenience wrapper for creating a simple number iterator
 */
public inline f<NumberIterator<Numeric>> range<Numeric>(Numeric begin, Numeric end) {
    return NumberIterator<Numeric>(begin, end);
}

/**
 * Convenience wrapper for creating a simple array iterator
 */
/*public inline f<ArrayIterator<I>> array<I>(I* array, unsigned long size) {
    return ArrayIterator<I>(array, size);
}*/