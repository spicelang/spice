// Imports
import "../ast/AstNodes" as ast;
import "../util/CodeLoc" as cl;

public type SemanticErrorType enum {
    REFERENCED_UNDEFINED_FUNCTION,
    REFERENCED_UNDEFINED_VARIABLE,
    REFERENCED_UNDEFINED_STRUCT,
    FUNCTION_AMBIGUITY,
    STRUCT_AMBIGUITY,
    VARIABLE_DECLARED_TWICE,
    FUNCTION_DECLARED_TWICE,
    GENERIC_TYPE_DECLARED_TWICE,
    STRUCT_DECLARED_TWICE,
    INTERFACE_DECLARED_TWICE,
    INTERFACE_METHOD_NOT_IMPLEMENTED,
    ENUM_DECLARED_TWICE,
    DUPLICATE_ENUM_ITEM_NAME,
    DUPLICATE_ENUM_ITEM_VALUE,
    GLOBAL_OF_TYPE_DYN,
    GLOBAL_OF_INVALID_TYPE,
    GLOBAL_CONST_WITHOUT_VALUE,
    MISSING_RETURN_STMT,
    INVALID_PARAM_ORDER,
    DTOR_MUST_BE_PROCEDURE,
    DTOR_WITH_PARAMS,
    OPERATOR_WRONG_DATA_TYPE,
    UNEXPECTED_DYN_TYPE,
    REASSIGN_CONST_VARIABLE,
    CONDITION_MUST_BE_BOOL,
    MISSING_MAIN_FUNCTION,
    FCT_PARAM_IS_TYPE_DYN,
    INVALID_BREAK_NUMBER,
    INVALID_CONTINUE_NUMBER,
    PRINTF_TYPE_ERROR,
    PRINTF_ARG_COUNT_ERROR,
    STD_NOT_FOUND,
    DUPLICATE_IMPORT_NAME,
    IMPORTED_FILE_NOT_EXISTING,
    CIRCULAR_DEPENDENCY,
    INVALID_MEMBER_ACCESS,
    SCOPE_ACCESS_ONLY_IMPORTS,
    UNKNOWN_DATATYPE,
    NUMBER_OF_FIELDS_NOT_MATCHING,
    FIELD_TYPE_NOT_MATCHING,
    ARRAY_SIZE_INVALID,
    ARRAY_INDEX_NOT_INT,
    ARRAY_ITEM_TYPE_NOT_MATCHING,
    EXPECTED_ARRAY_TYPE,
    SIZEOF_DYNAMIC_SIZED_ARRAY,
    RETURN_WITHOUT_VALUE_RESULT,
    RETURN_WITH_VALUE_IN_PROCEDURE,
    DYN_POINTERS_NOT_ALLOWED,
    DYN_ARRAYS_NOT_ALLOWED,
    GENERIC_TYPE_NOT_IN_TEMPLATE,
    SPECIFIER_AT_ILLEGAL_CONTEXT,
    INSUFFICIENT_VISIBILITY,
    TID_INVALID,
    JOIN_ARG_MUST_BE_TID,
    EXPECTED_GENERIC_TYPE,
    EXPECTED_STRUCT_TYPE,
    EXPECTED_INTERFACE_TYPE,
    INTERFACE_WITH_TEMPLATE_LIST,
    EXPECTED_VALUE,
    EXPECTED_TYPE,
    UNSAFE_OPERATION_IN_SAFE_CONTEXT,
    ASSERTION_CONDITION_BOOL,
    ARRAY_INDEX_OUT_OF_BOUNDS,
    RESERVED_KEYWORD,
    COMING_SOON_SA
}

public type SemanticError struct {
    string message
}

public p SemanticError.ctor(const ast::AstNode* node, const SemanticErrorType errorType, const string message) {
    this.errorMessage = "[Error|Semantic] " + node.codeLoc.toPrettyString() + ":\n" + this.getMessagePrefix(errorType) +
            ": " + message + "\n\n" + node.errorMessage;
}

/**
 * Get the prefix of the error message for a particular error
 *
 * @param type Type of the error
 * @return Prefix string for the error type
 */
f<string> SemanticError.getMessagePrefix(const SemanticErrorType errorType) {
    if errorType == SemanticErrorType.REFERENCED_UNDEFINED_FUNCTION { return "Referenced undefined function"; }
    if errorType == SemanticErrorType.REFERENCED_UNDEFINED_VARIABLE { return "Referenced undefined variable"; }
    if errorType == SemanticErrorType.REFERENCED_UNDEFINED_STRUCT { return "Referenced undefined struct"; }
    if errorType == SemanticErrorType.FUNCTION_AMBIGUITY { return "Function ambiguity"; }
    if errorType == SemanticErrorType.STRUCT_AMBIGUITY { return "Struct ambiguity"; }
    if errorType == SemanticErrorType.VARIABLE_DECLARED_TWICE { return "Multiple declarations of the same variable"; }
    if errorType == SemanticErrorType.FUNCTION_DECLARED_TWICE { return "Multiple declarations of a function/procedure"; }
    // ToDo: Extend
    return "Unknown error";
}