type Person struct {
    string* firstName
    string* lastName
    int age
}

type Person struct {
    int age
    double* height
    Person* person
}

f<int> main() {}