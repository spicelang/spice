#[test]
f<bool> testAdd() {
    return false; // Returning false means the test failed
}
