import "std/os/thread-pool";
import "std/time/delay";

f<int> main() {
    ThreadPool tp = ThreadPool(3s);
    tp.enqueue(p() [[async]] {
        delay(50);
        printf("Hello from task 1\n");
    });
    tp.enqueue(p() [[async]] {
        delay(100);
        printf("Hello from task 2\n");
    });
    tp.enqueue(p() [[async]] {
        delay(150);
        printf("Hello from task 3\n");
    });
    tp.enqueue(p() [[async]] {
        delay(200);
        printf("Hello from task 4\n");
    });
    tp.enqueue(p() [[async]] {
        delay(250);
        printf("Hello from task 5\n");
    });
    tp.enqueue(p() [[async]] {
        delay(300);
        printf("Hello from task 6\n");
    });
    tp.enqueue(p() [[async]] {
        delay(350);
        printf("Hello from task 7\n");
    });
    tp.enqueue(p() [[async]] {
        delay(400);
        printf("Hello from task 8\n");
    });
    tp.enqueue(p() [[async]] {
        delay(450);
        printf("Hello from task 9\n");
    });
    tp.enqueue(p() [[async]] {
        delay(500);
        printf("Hello from task 10\n");
    });
    tp.start();
    tp.join();
}

/*import "std/os/thread-pool";

f<int> main() {
    int testVar = 123;
    ThreadPool tp = ThreadPool(3s);
    dyn proc = p() [[async]] {
        printf("Hello from inside: %d\n", testVar);
    };
    tp.enqueue(proc);
    tp.start();
    tp.join();
    printf("TestVar: %d\n", testVar);
}*/

/*f<int> main() {
    int i = 123; // Captured by ref
    int j = 321; // Captured by val
    dyn lambda = p() {
        printf("Hello from inside: %d\n", i);
        i++;
        i += j;
        printf("Hello from inside: %d\n", i);
    };
    lambda();
    printf("Hello from outside: %d\n", i);
}*/

/*type Visitable interface {
    p print();
}

type Test1 struct : Visitable {
    int f1
}

p Test1.print() {
    printf("Foo: %d", this.f1);
}

f<int> main() {
    Test1 t1 = Test1{123};
    Visitable* v = &t1;
    v.print();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";

f<int> main() {
    Lexer lexer = Lexer("./file.spice");
    Parser parser = Parser(lexer);
    parser.parse();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "std/time/timer";

f<int> main() {
    Timer timer = Timer();
    timer.start();
    Lexer lexer = Lexer("./file.spice");
    unsigned long i = 1l;
    while (!lexer.isEOF()) {
        Token token = lexer.getToken();
        //printf("Token %d: ", i);
        //token.print();
        lexer.advance();
        i++;
    }
    timer.stop();
    printf("Tokens: %d, Time: %d\n", i, timer.getDurationInMillis());
}*/