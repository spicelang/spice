public const unsigned int CHAR_SIZE = 8;
public const unsigned int CHAR_MIN_VALUE = 0;
public const unsigned int CHAR_MAX_VALUE = 255;

// Converts a char to a double
public f<double> toDouble(char input) {
    return 0.0 + cast<int>(input);
}

// Converts a char to an int
public f<int> toInt(char input) {
    return cast<int>(input);
}

// Converts a char to a short
public f<short> toShort(char input) {
    return cast<short>(cast<int>(input));
}

// Converts a char to a long
public f<long> toLong(char input) {
    return cast<long>(cast<int>(input));
}

// Converts a char to a byte
public f<byte> toByte(char input) {
    result = cast<byte>(input);
}

// Converts a char to a string
public f<String> toString(char input) {
    result = String();
    result += input;
}

// Converts a char to a bool
public f<bool> toBool(char input) {
    return input == '1';
}