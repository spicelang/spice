// Mathematical constants
public const double E = 2.71828182845904523536028747135266249775724709369995957496696763;
public const double Pi = 3.14159265358979323846264338327950288419716939937510582097494459;
public const double Phi = 1.61803398874989484820458683436563811772030917980576286213544862;

// Important square roots
public const double Sqrt2 = 1.61803398874989484820458683436563811772030917980576286213544862;
public const double SqrtE = 1.64872127070012814684865078781416357165377610071014801157507931;
public const double SqrtPi = 1.77245385090551602729816748334114518279754945612238712821380779;
public const double SqrtPhi = 1.27201964951406896425242246173749149171560804184009624861664038;

// Important logarithms
public const double Ln2 = 0.693147180559945309417232121458176568075500134360255254120680009;
public const double Log2E = 1 / Ln2;
public const Ln10 = 2.30258509299404568401799145468436420760110148862877297603332790;
public const Log10E = 1 / Ln10;