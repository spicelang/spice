public const int SIZE = 32;
public const int MIN_VALUE = -2147483648;
public const int MAX_VALUE = 2147483647;

// Converts an int to a double
public f<double> toDouble(int input) {
    return 0.0 + input;
}

// Converts an int to a short
public f<short> toShort(int input) {
    return (short) input;
}

// Converts an int to a long
public f<long> toLong(int input) {
    return (long) input;
}

// Converts an int to a byte
public f<byte> toByte(int input) {
    return (byte) input;
}

// Converts an int to a char
public f<char> toChar(int input) {
    return (char) input;
}

// Converts an int to a string
public f<string> toString(const int input) {
    if input == 0 { return "0"; }

    string str;
    bool isNeg = input < 0;
    unsigned int uInput = isNeg ? -input : input;

    while (uInput != 0) {
        str.append((char) (uInput % 10 + 48 /* ASCII for '0' */));
        uInput = uInput / 10;
    }
    if isNeg { str.append('-'); }

    //return str.reverse();
    return str;
}

// Converts an int to a boolean
public f<bool> toBool(int input) {
    return input >= 1;
}

// Check if the input is a power of two
public f<bool> isPowerOfTwo(int input) {
    return (input & (input - 1)) == 0;
}