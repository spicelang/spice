public type ThreadFactory struct {
    unsigned long nextSuffix
}

public p ThreadFactory.ctor() {
    this.nextSuffix = 0l;
}

public f<int> ThreadFactory.getNextFunctionSuffix() {
    return this.nextSuffix++;
}

public f<bool> ThreadFactory.isUsingThreads() {
    return this.nextSuffix > 0l;
}