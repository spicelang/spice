f<int> main() {
    printf("Hi.\n");
}

1