ext f<byte*> malloc(int);

f<int> test(string input) {
    return 12;
}

p invoke(f<int>(string) fctPtr) {
    fctPtr("string");
}

f<int> main() {
    f<int>(string) testFct = test;
    invoke(testFct);
}