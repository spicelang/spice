type Test struct {
    int i = 12
    string s = "test"
}

f<int> main() {
    Test t;
    printf("Int: %d\n", t.i);
    printf("String: %s\n", t.s);
}

/*type TestStruct struct {
    int a = 123
    short b = 1s
}

f<int> main() {
    TestStruct ts;
    printf("%d %d\n", ts.a, ts.b);
}*/