// Link WinSock library
#![core.linux.linker.flag = "-lws2_32"]

// Import common logic
import "std/net/socket";

// Type defs
type SAFamilyT alias unsigned short;

// Constants
const unsigned short REQUESTED_WSA_VERSION = 514s;

type WSAData struct {
    unsigned short wVersion
    unsigned short wHighVersion
    unsigned short iMaxSockets
    unsigned short iMaxUdpDg
    char* lpVendorInfo
    char[257] szDescription
    char[129] szSystemStatus
}

// External functions
ext f<int> WSAStartup(short, WSAData*);
ext f<int> WSACleanup();
ext f<int> socket(int /*sockfd*/, int /*type*/, int /*protocol*/);
ext f<int> bind(int /*sockfd*/, SockAddrIn* /*address*/, SockLenT /*address_len*/);
ext f<int> listen(int /*sockfd*/, int /*backlog*/);
ext f<int> accept(int /*sockfd*/, SockAddrIn*, SockLenT /*address_len*/);
ext f<int> close(int /*sockfd*/);
ext f<unsigned int> htonl(unsigned int /*hostlong*/);      // Fairly simple to re-implement in Spice
ext f<unsigned short> htons(unsigned short /*hostshort*/); // Fairly simple to re-implement in Spice

type SockAddr struct {
    SAFamilyT saFamily // Address family
    char[] saData      // Socket address
}

type SockAddrStorage struct {
    SAFamilyT ssFamily // Address family
}

// Represents an IPv4 address
public type InAddr struct {
    InAddrT addr
}

// Represents an IPv6 address
public type In6Addr struct {
    unsigned byte[16] addr
}

public type SockAddrIn struct {
    unsigned short sinFamily // AF_INET
    InPortT sinPort          // Port number
    InAddr sinAddr           // IPv4 address
}

public type SockAddrIn6 struct {
    unsigned short sin6Family // AF_INET6
    InPortT sin6Port          // Port number
    unsigned int sin6FlowInfo // IPv6 flow info
    In6Addr sin6Addr          // IPv6 address
    unsigned int sin6ScopeId  // Set of interfaces for a scope
}

public type SockAddrUn struct {

}

public type Socket struct {
    int sockFd // Actual socket
    int connFd // Current connection
}

/**
 * Accept an incoming connection to the socket and save the connection file desceiptor
 * to the socket object.
 *
 * @return Connection file descriptor
 */
public f<Result<int>> Socket.acceptConnection() {
    SockAddrIn cliAddr = SockAddrIn {};
    this.connFd = accept(this.sockFd, &cliAddr, 16u /* hardcoded sizeof(cliAddr) */);
    if this.connFd == -1 { return err<int>(Error("Error while accepting connection")); }
    return ok(this.connFd);
}

/**
 * Closes the socket. This method should always be called by the user before exiting the program.
 *
 * @return Closing the connection was successful or not
 */
public f<bool> Socket.close() {
    return close(this.sockFd) == 0 && WSACleanup() == 0;
}

/**
 * Opens a TCP server socket and exposes it to the given port.
 * The maxWaitingConnections defines the maximum length to which the queue of pending connections may grow. If a
 * connection request arrives when the queue is full, the client may receive an error with an indication of
 * ECONNREFUSED or, if the underlying protocol support retransmission, the request may be ignored so that a later
 * reattempt at connection succeeds.
 *
 * @param port Port to open the socket on
 * @param maxWaitingConnections Maximum size of the queue of pending client connections
 * @return Socket file descriptor
 */
public f<Result<Socket>> openServerSocket(unsigned short port, int maxWaitingConnections = 5) {
    // Initialize WSA
    WSAData wsaData = WSAData{};
    if WSAStartup(REQUESTED_WSA_VERSION, &wsaData) != 0 { return err<Socket>(Error("Error initializing WSA")); }

    // Create socket file descriptor
    const int sockFd = socket(AF_INET, SOCK_STREAM, IPPROTO_IP);
    if sockFd == -1 { return err<Socket>(Error("Error creating socket")); }

    // Construct socket object
    const Socket s = Socket { sockFd, /*connFd*/ 0 };
    SockAddrIn servAddr = SockAddrIn { cast<short>(AF_INET), htons(port), InAddr { INADDR_ANY }};

    // Bind to target address
    int bindResult = bind(sockFd, &servAddr, 16u /* hardcoded sizeof(servaddr) */);
    if bindResult != 0 { return err<Socket>(Error("Error binding to address")); }

    // Start listening for incoming connections
    int listenResult = listen(s.sockFd, maxWaitingConnections);
    if listenResult != 0 { return err<Socket>(Error("Error listening on address")); }

    return ok(s);
}
