f<int> main() {
    f<int>(int, int) add = f<int>(int x, int y) {
        return "String";
    };
}