f<int> main() {
    string output = "Hello world!";
    sout.println(output);
}