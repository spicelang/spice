public type NestedSocket struct {
    public string testString
    long _testLong
}

public type Socket struct {
    public int sock // Actual socket
    short _errorCode
    public NestedSocket nested
}

public f<Socket> openServerSocket(unsigned short _port) {
    dyn nested = NestedSocket { "Test", 2345l };
    return Socket{ 2, 0s, nested };
}