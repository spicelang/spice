f<int> main() {
    f<int>(int, int) add = f<dyn>(int x, int y) {
        return x + y;
    };
}