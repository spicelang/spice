import "std/type/bool" as boolTy;

f<int> main() {
    printf("Result: %d", boolTy.toInt(true));
}