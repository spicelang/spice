f<int> main() {
    string s;
    len(s);
}