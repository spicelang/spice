public type Vector1 struct {
    public int i2
}

public type Vector struct {
    public Vector1 i1
}

public p Vector1.ctor() {

}