f<bool> functionTrue() {
    printf("Function True\n");
    return true;
}

f<bool> functionFalse() {
    printf("Function False\n");
    return false;
}

f<int> main() {
    // Short circuiting for logical and op
    printf("Logical and evaluated to: %d\n", functionFalse() && functionTrue());

    // Short circuiting for logical or op
    printf("Logical or evaluated to: %d\n", functionTrue() || functionFalse());
}

/*type T string|char;

type TestStruct<T> struct {
    T base
    int test
}

f<int> main() {
    TestStruct<char> s = TestStruct<char>{ 'a', 1 };
    s.printTest();
}

p TestStruct.printTest() {
    printf("Test: %d\n", this.getTest());
}

f<int> TestStruct.getTest() {
    if this.test == 1 {
        this.test++;
        this.printTest();
    }
    return this.test;
}*/

/*ext<byte*> malloc(long);
ext free(byte*);

f<int> main() {
    byte* address = malloc(1l);
    *address = (byte) 12;
    free(address);
}*/

/*f<int> main() {
    int[10] a;
    for int i = 0; i < len(a); i++ {
        a[i] = 1;
    }
    printf("Cell [3]: %d", a[3]);
}*/