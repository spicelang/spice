f<int> main() {
    char* s = "abc";
    printf("%s\n", (char*) s);
}