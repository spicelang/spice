f<int> main() {
    long l = 1234l;
    long* lPtr = &l;
    int* iPtr = (int*) lPtr;
    printf("Int: %d\n", *iPtr);
}