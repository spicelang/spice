f<int> main() {
    // Plus
    printf("Result: %s\n", String("Hello ") + String("World!"));
    String s1 = String("Hello ") + String("World!");
    printf("Result: %s\n", s1);
    printf("Result: %s\n", s1 + " Hi!");
    printf("Result: %s\n", String("Hi! ") + s1);
    printf("Result: %s\n", s1 + s1);
    printf("Result: %s\n", s1 + " " + s1);
    printf("Result: %s\n", String("Prefix ") + s1 + " Suffix");

    // Mul
    printf("Result: %s\n", 4s * String("Hi"));
    String s2 = String("Hello ") * 5;
    printf("Result: %s\n", s2);
    printf("Result: %s\n", 20 * String('a'));
    String s3 = 2 * String('c') * 7;
    printf("Result: %s\n", s3);
    printf("Result: %s\n", String("One") * 1);

    // Equals raw
    printf("Equal raw: %d\n", "Hello World!" == "Hello Programmers!");
    printf("Equal raw: %d\n", "Hello" == "Hell2");
    printf("Equal raw: %d\n", "Hello" == "Hello");

    // Equals
    printf("Equal: %d\n", String("Hello World!") == String("Hello Programmers!"));
    printf("Equal: %d\n", String("Hello") == String("Hell2"));
    printf("Equal: %d\n", String("Hello") == String("Hello"));

    // Not equals raw
    printf("Non-equal raw: %d\n", "Hello World!" != "Hello Programmers!");
    printf("Non-equal raw: %d\n", "Hello" != "Hell2");
    printf("Non-equal raw: %d\n", "Hello" != "Hello");

    // Not equals
    printf("Non-equal: %d\n", String("Hello World!") != String("Hello Programmers!"));
    printf("Non-equal: %d\n", String("Hello") != String("Hell2"));
    printf("Non-equal: %d\n", String("Hello") != String("Hello"));

    // PlusEquals
    String s4 = String("Hello");
    s4 += 'l';
    printf("Result: %s\n", s4);
    String s5 = String("Hi");
    s5 += " World!";
    printf("Result: %s\n", s5);

    // MulEquals
    String s6 = String("Hi");
    s6 *= 3;
    printf("Result: %s\n", s6);
}

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";
import "../../src-bootstrap/ast/ast-nodes";

f<int> main() {
    Lexer lexer = Lexer("./test-file.spice");
    Parser parser = Parser(lexer);
    ASTEntryNode* entryNode = parser.parse();
}*/

/*f<int> main() {
    int i = 123; // Captured by ref
    int j = 321; // Captured by val
    dyn lambda = p() {
        printf("Hello from inside: %d\n", i);
        i++;
        i += j;
        printf("Hello from inside: %d\n", i);
    };
    lambda();
    printf("Hello from outside: %d\n", i);
}*/

/*type Visitable interface {
    p print();
}

type Test1 struct : Visitable {
    int f1
}

p Test1.print() {
    printf("Foo: %d", this.f1);
}

f<int> main() {
    Test1 t1 = Test1{123};
    Visitable* v = &t1;
    v.print();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";

f<int> main() {
    Lexer lexer = Lexer("./file.spice");
    Parser parser = Parser(lexer);
    parser.parse();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "std/time/timer";

f<int> main() {
    Timer timer = Timer();
    timer.start();
    Lexer lexer = Lexer("./file.spice");
    unsigned long i = 1l;
    while (!lexer.isEOF()) {
        Token token = lexer.getToken();
        //printf("Token %d: ", i);
        //token.print();
        lexer.advance();
        i++;
    }
    timer.stop();
    printf("Tokens: %d, Time: %d\n", i, timer.getDurationInMillis());
}*/