f<int> main() {
    int[3] a = [1, 2, 3];
    int* aPtr = a;
    printf("%d\n", *aPtr);
    unsafe {
        aPtr++;
    }
    printf("%d\n", *aPtr);
}

/*import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

f<int> main() {
    DefaultMemoryManager defaultMemoryManager;
    IMemoryManager* memoryManager = &defaultMemoryManager;
    BlockAllocator<int> allocator = BlockAllocator<int>(memoryManager, 10l);
}*/