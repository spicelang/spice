

public type QualType struct {

}