f<int> main() {
    int arraySize = 4;
    int[arraySize] intArray;
    intArray[0] = 10;
    intArray[1] = 12;
    intArray[2] = 7;
    printf("Test: %d\n", intArray[0]);
    printf("Size: %d\n", len(intArray));
}