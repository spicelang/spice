f<int> main() {
    String s = String("Dies ist ein Test. Und weil das ein Test ist, ist es ein Test.");
    long replaced = s.replaceAll("ist", "wart");
    printf("Result: %d\n", replaced);
    printf("Result: %s\n", s.getRaw());
}