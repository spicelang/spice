// Std imports
import "std/type/any";

public type IAbstractAstVisitor interface {
    f<Any> visitEntry(ASTEntryNode*);
    f<Any> visitMainFctDef(ASTMainFctDefNode*);
    f<Any> visitFctDef(ASTFctDefNode*);
    f<Any> visitProcDef(ASTProcDefNode*);
}