import "std/os/syscall";

f<int> main() {
    // Use write syscall to print "Hello syscall!"
    const string str = "Hello syscall!";
    syscall(SYSCALL_WRITE, /*fd = stdout*/ 1, /* buffer */ str, len(str));
}