ext f<unsigned int> snprintf(char*, unsigned long, string, ...);

f<int> main() {

}