//import "std/os/thread";

ext f<int> pthread_create(byte* /*thread*/, byte* /*attr*/, p() /*start_routine*/, byte* /*arg*/);

type EmptyParams struct {}

p threadRoutine() {
    //printf("Hello from thread: %p\n", getThreadId());
    printf("Test");
}

f<int> main() {
    byte tid;
    EmptyParams emptyParams;
    unsafe {
        pthread_create(&tid, nil<byte*>, threadRoutine, (byte*) &emptyParams);
    }

    //Thread t1 = Thread();
    //Thread t2 = Thread(threadRoutine);
    //t1.join();
    //t2.join();
}