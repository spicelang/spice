// Std imports
import "std/text/stringstream";

// Own imports
import "bootstrap/reader/code-loc";

public type CliErrorType enum {
    INCOMPLETE_TARGET_TRIPLE,
    INVALID_TARGET_TRIPLE,
    SOURCE_FILE_MISSING,
    INCOMPATIBLE_OPTIONS,
    NON_ZERO_EXIT_CODE,
    FEATURE_NOT_SUPPORTED_FOR_TARGET,
    FEATURE_NOT_SUPPORTED_WHEN_DOCKERIZED,
    INVALID_BUILD_MODE,
    INVALID_OUTPUT_CONTAINER,
    INVALID_SANITIZER
}

/**
 * Custom exception for errors, occurring when linking the output executable
 */
public type CliError struct {
    String errorMessage
}

/**
 * @param errorType Type of the error
 * @param message Error message suffix
 */
public p CliError.ctor(const CliErrorType errorType, const string message) {
    StringStream msg;
    msg << "[Error|CLI] " << this.getMessagePrefix(errorType) << ": " << message;
    this.errorMessage = msg.str();
}

/**
 * Get the prefix of the error message for a particular error
 *
 * @param errorType Type of the error
 * @return Prefix string for the error type
 */
f<string> CliError.getMessagePrefix(const CliErrorType errorType) {
    switch errorType {
        case CliErrorType::INCOMPLETE_TARGET_TRIPLE: { return "Incomplete target triple"; }
        case CliErrorType::INVALID_TARGET_TRIPLE: { return "Invalid target triple"; }
        case CliErrorType::SOURCE_FILE_MISSING: { return "Source file missing"; }
        case CliErrorType::INCOMPATIBLE_OPTIONS: { return "Incompatible options"; }
        case CliErrorType::NON_ZERO_EXIT_CODE: { return "Non-zero exit code"; }
        case CliErrorType::FEATURE_NOT_SUPPORTED_FOR_TARGET: { return "Feature is not supported for this target"; }
        case CliErrorType::FEATURE_NOT_SUPPORTED_WHEN_DOCKERIZED: { return "Feature not supported when dockerized"; }
        case CliErrorType::INVALID_BUILD_MODE: { return "Invalid build mode"; }
        case CliErrorType::INVALID_OUTPUT_CONTAINER: { return "Invalid output container"; }
        case CliErrorType::INVALID_SANITIZER: { return "Invalid sanitizer"; }
        default: { panic(Error("Unknown error")); }
    }
}