f<int> main() {
    int test = "Test";
}