import "bootstrap/util/system-util";

f<int> main() {
    printf("GCC installed: %s\n", isCommandAvailable("gcc") ? "yes" : "no");
    printf("Graphviz installed: %s\n", isGraphvizInstalled() ? "yes" : "no");
    ExternalBinaryFinderResult linkerInvoker = findLinkerInvoker();
    assert linkerInvoker.path.contains("clang") || linkerInvoker.path.contains("gcc");
    printf("All assertions passed!");
}