f<int> main(int argc, string[] argv) {
    printf("Argc: %d\n", argc);
    printf("Argv no. 0: %s\n", argv[0]);
    if (argc > 1) {
        printf("Argv no. 1: %s\n", argv[1]);
    }
}