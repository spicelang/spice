import "std/iterators/iterable";

// Generic type definitions
type T int|long|short;

/**
 * A NumberIterator in Spice can be used to iterate over a range of numbers
 */
public type NumberIterator<T> struct : Iterable<T> {
    T lowerBound // Inclusive
    T upperBound // Inclusive
    unsigned long cursor
}

public p NumberIterator.ctor(T lowerBound, T upperBound) {
    this.lowerBound = lowerBound;
    this.upperBound = upperBound;
    this.cursor = 0l;
}

/**
 * Check if the number range has another number
 *
 * @return true or false
 */
public inline const f<bool> NumberIterator.hasNext() {
    return this.lowerBound + this.cursor <= this.upperBound;
}

/**
 * Returns the current number of the number range and moves the cursor to the next item
 *
 * @return current item
 */
public inline f<T> NumberIterator.next() {
    assert this.hasNext();
    T currentItem = this.get();
    this.cursor++;
    return currentItem;
}

/**
 * Returns the current number of the number range
 */
public inline f<T> NumberIterator.get() {
    return (T) (this.lowerBound + this.cursor);
}