// Std imports
import "std/data/vector";

// Own imports
import "bootstrap/symboltablebuilder/qual-type-intf";
import "bootstrap/symboltablebuilder/type";
import "bootstrap/symboltablebuilder/type-chain";
import "bootstrap/symboltablebuilder/type-qualifiers";

public type QualType struct : IQualType {
    const Type* rawType
    TypeQualifiers qualifiers
}

public p QualType.ctor(SuperType superType) {

}

public p QualType.ctor(SuperType superType, const String& subType) {

}

public p QualType.ctor(const Type* rawType, TypeQualifiers qualifiers) {
    this.rawType = rawType;
    this.qualifiers = qualifiers;
}

public type QualTypeList alias Vector<QualType>;