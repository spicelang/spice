// Std imports
import "std/text/stringstream";

// Own imports
import "bootstrap/util/code-loc";

public type LinkerErrorType enum {
    LINKER_NOT_FOUND,
    LINKER_ERROR
}

/**
 * Custom exception for errors, occurring when linking the output executable
 */
public type LinkerError struct {
    string errorMessage
}

/**
 * @param type Type of the error
 * @param message Error message suffix
 */
public p LinkerError.ctor(const LinkerErrorType errorType, const string message) {
    StringStream msg;
    msg << "[Error|Linker] " << this.getMessagePrefix(errorType) << ": " << message;
    this.errorMessage = msg.str();
}

/**
 * Get the prefix of the error message for a particular error
 *
 * @param errorType Type of the error
 * @return Prefix string for the error type
 */
f<string> LinkerError.getMessagePrefix(const LinkerErrorType errorType) {
    switch errorType {
        case LinkerErrorType::LINKER_NOT_FOUND: { return "Linker not found"; }
        case LinkerErrorType::LINKER_ERROR: { return "Linker error occurred"; }
        default: { panic(Error("Unknown error")); }
    }
}