// Imports

public type SymbolTableEntry struct {

}

public p SymbolTableEntry.ctor() {

}