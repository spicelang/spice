import "std/type/long" as longTy;

f<int> main() {
    // toDouble()
    double asDouble = longTy.toDouble(123l);
    assert asDouble == 123.0;

    // toInt()
    int asInt = longTy.toInt(459873l);
    assert asInt == 459873;

    // toShort()
    short asShort = longTy.toShort(-345l);
    assert asShort == -345s;

    // toByte()
    byte asByte = longTy.toByte(12l);
    assert asByte == (byte) 12;

    // toChar()
    char asChar = longTy.toChar(66l);
    assert asChar == 'B';

    // toString()
    //string asString = longTy.toString(12345l);
    //assert asString == "12345";
    //printf("Str: %s\n", asString);

    // toBool()
    bool asBool1 = longTy.toBool(1l);
    assert asBool1 == true;
    bool asBool2 = longTy.toBool(0l);
    assert asBool2 == false;

    // isPowerOfTwo()
    assert longTy.isPowerOfTwo(16l);
    assert !longTy.isPowerOfTwo(31l);

    printf("All assertions succeeded");
}