type A dyn;

public p printFormat<A>(A element) {
    printf("Test");
    /*printf("Sizeof output: %d\n", sizeof(element));*/
}