import "std/time/delay" as delay;
import "std/os/cpu" as cpu;

type Mutex struct {
	bool occupied
}

p Mutex.acquire() {
	while this.occupied {
		cpu.yield();
	}
	this.occupied = true;
}

p Mutex.abandon() {
	this.occupied = false;
}