// Imports
import "std/io/cli-parser";

import "SourceFile";
import "CliInterface";
import "global/GlobalResourceManager";

/**
 * Compile main source file. All files, that are included by the main source file will be resolved recursively.
 *
 * @param options Command line options
 */
f<int> compileProject(const CliOptions& options) {
    // Instantiate GlobalResourceManager
    dyn resourceManager = GlobalResourceManager(options);

    // Create source file instance for main source file
    dyn mainSourceFile = SourceFile(options, nil<SourceFile*>, "root", options.mainSourceFile, false);

    // Run compile pipeline for main source file. All dependent source files are triggered by their parents
    mainSourceFile.runFrontEnd();
    mainSourceFile.runMiddleEnd();
    mainSourceFile.runBackEnd();

    // Link the target executable (link object files to executable)
    if !options.execute {
        resourceManager.linker.prepare();
        resourceManager.linker.link();
    }

    // Print compiler warnings
    mainSourceFile.collectAndPrintWarnings();

    if options.execute {
        return mainSourceFile.execute();
    }

    return 0;
}

/**
 * Entry point to the Spice compiler
 *
 * @param argc Argument count
 * @param argv Argument vector
 * @return Return code
 */
f<int> main(int argc, string[] argv) {
    // Initialize command line parser
    CliInterface cli;
    cli.createInterface();
    if (cli.parse(argc, argv) != 0) {
        return 1;
    }
    if (!cli.shouldCompile) {
        return 0;
    }
    cli.enrich();   // Prepare the cli options

    // Kick off the compiling process
    return compileProject(cli.cliOptions);
}