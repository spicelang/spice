f<int> main() {
    dyn test;
}