import "std/data/vector" as v;

f<int> main() {
    dyn vec = v.Vector<int>();
    vec.pushBack(12);

}