import "std/os/os";
import "std/data/vector";
import "std/io/filepath";

// Generic types
type T bool|string|String|int|long|short|FilePath;

// Enums
type CliOptionMode enum { SET_VALUE, CALL_CALLBACK }

public type CliOption<T> struct {
    String name
    String description
    Vector<String> aliases
    CliOptionMode mode
    T& targetVariable
    p(T&) callback
}

public p CliOption.ctor(const String& name, T& targetVariable, const String& description) {
    this.name = name;
    this.description = description;
    this.mode = CliOptionMode::SET_VALUE;
    this.targetVariable = targetVariable;
}

public p CliOption.ctor(const String& name, p(T&) callback, const String& description) {
    this.name = name;
    this.description = description;
    this.mode = CliOptionMode::CALL_CALLBACK;
    this.callback = callback;
}

public const f<const String&> CliOption.getName() {
    return this.name;
}

public const f<const String&> CliOption.getDescription() {
    return this.description;
}

public p CliOption.addAlias(string optionName) {
    this.aliases.pushBack(String(optionName));
}

public p CliOption.addAlias(const String& optionName) {
    this.aliases.pushBack(optionName);
}

public const f<const Vector<String>&> CliOption.getAliases() {
    return this.aliases;
}

public p CliOption.setTargetValue(T value) {
    if this.mode == CliOptionMode::SET_VALUE {
        this.targetVariable = value;
    }
}

public p CliOption.callCallback(T& value) {
    if this.mode == CliOptionMode::CALL_CALLBACK {
        p(T&) cb = this.callback;
        cb(value);
    }
}