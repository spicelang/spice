public type TestAlias alias int;