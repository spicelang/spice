f<int> main() {
    assert true;
    printf("First assertion was true\n");

    assert 1 != 1;
    printf("Unreachable");
}