/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

f<int> main() {
    int[10] intArray = { 1, 2, 4, 8, 16, 32, 64, 128, 256, 512, 1024 };
    printf("intArray[3]: %d\n", intArray[3]);
    printf("intArray[7]: %d\n", intArray[7]);
    printf("intArray[9]: %d\n", intArray[9]);
}