f<int> main() {
    return 1-2;
}