f<int> main() {
    String s1 = String("Hello World!");
    printf("S1: %s\n", s1);
    String s2 = String(s1);
    s2 += " Hi!";
    printf("S1: %s\n", s1);
    printf("S2: %s\n", s2);
}

/*type TestStruct struct {
    long test
}

f<TestStruct&> operator++(TestStruct& ts) {
    ts.test++;
    return ts;
}

f<int> main() {
    TestStruct ts = TestStruct{ 123l };
    TestStruct& output = ts++;
    ts.test++;
    assert output.test == 125l;
    assert ts.test == 125l;
}*/