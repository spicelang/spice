f<int> main() {
    double calcResult = 1 != 2 ? false : 1.0;
}