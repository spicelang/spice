// Std imports
import "std/io/filepath";
import "std/io/file";
import "std/type/result";
import "std/type/error";

// Own import
import "../reader/code-loc";

public type Reader struct {
    File file
    string filename
    char curChar = '\0'
    unsigned long line = 1l
    unsigned long col = 0l
}

public p Reader.ctor(const string inputFileName) {
    this.filename = inputFileName;
    Result<File> result = openFile(inputFileName, MODE_READ);
    if !result.isOk() {
        panic(Error("Source file cannot be opened"));
    }
    this.file = result.unwrap();
}

public p Reader.dtor() {
    this.file.close();
}

/**
 * @brief Get the previously read character
 *
 * @return char Last character
 */
public f<char> Reader.getChar() {
    return this.curChar;
}

/**
 * @brief Get the code location of the previously read character
 *
 * @return CodeLoc Code location
 */
public f<CodeLoc> Reader.getCodeLoc() {
    return CodeLoc(this.line, this.col, this.filename);
}

/**
 * @brief Advance the reader by one character
 */
public p Reader.advance() {
    assert !this.isEOF();
    this.curChar = (char) this.file.readChar();
    if this.curChar == '\n' {
        this.line++;
        this.col = 0l;
    }
    this.col++;
}

/**
 * @brief Advance the reader by one character and check if this char equals the
 * expected
 *
 * @param c Expected char
 */
public p Reader.expect(char c) {
    assert this.curChar == c;
    this.advance();
}

/**
 * @brief Check if we are at the end of the input file
 *
 * @return At the end or not
 */
public f<bool> Reader.isEOF() {
    return this.file.isEOF();
}