public type IInterface interface {

}
