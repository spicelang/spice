public type Test struct {
    public int t
}

public p Test.ctor() {

}

//const int globalTestVar = 123;