// Imports
import "std/math/const";
import "std/type/double" as doubleType;

// Generic type defs
type Numeric double|int|short|long;
type WholeNumber int|short|long;

/**
 * Calculate absolute value of the input
 *
 * @param input Input number
 * @return Absulute value of input
 */
public inline f<Numeric> abs<Numeric>(Numeric input) {
    return input < 0 ? -input : input;
}

/**
 * Calculate the maximum of two inputs
 *
 * @param input1 First input
 * @param input2 Second input
 * @return Maximum of inputs
 */
public inline f<Numeric> max<Numeric>(Numeric input1, Numeric input2) {
    return input1 > input2 ? input1 : input2;
}

/**
 * Calculate the minimum of two inputs
 *
* @param input1 First input
* @param input2 Second input
* @return Minimum of inputs
 */
public inline f<Numeric> min<Numeric>(Numeric input1, Numeric input2) {
    return input1 < input2 ? input1 : input2;
}

/**
 * Truncate the number to a whole number
 *
 * @param input Intput number
 * @return Rounding result
 */
public inline f<int> trunc(double input) {
    return doubleType::toInt(input);
}

/**
 * Round the input number down
 *
 * @param input Intput number
 * @return Rounding result
 */
public inline f<int> floor(double input) {
    const int truncated = trunc(input);
    if input >= 0.0 { return truncated; }
    return truncated == input ? truncated : truncated - 1;
}

/**
 * Round the input number up
 *
 * @param input Intput number
 * @return Rounding result
 */
public inline f<int> ceil(double input) {
    const int truncated = trunc(input);
    if input <= 0.0 { return truncated; }
    return truncated == input ? truncated : truncated + 1;
}

/**
 * Round the input number to a whole number
 * Note: 0.499999 is rounded down to 0, 0.5 is rounded up to 1.
 *
 * @param input Input number
 * @return Rounding result
 */
public inline f<int> round(double input) {
    return cast<int>(input + (input >= 0.0 ? 0.5 : -0.5));
}

/**
 * Round the input number to the given number of decimal places
 * Note: For 2 places 0.444 is rounded down to 0.44, 0.445 is rounded up to 0.45.
 *
 * @param input Input number
 * @param places Number of decimal places
 * @param Rounding result
 */
public inline f<double> round(double input, unsigned int places) {
    double factor = 1.0;
    for unsigned int i = 0u; i < places; i++ {
        factor *= 10.0;
    }
    return cast<int>(input * factor + (input >= 0.0 ? 0.5 : -0.5)) / factor;
}

/**
 * Convert degrees to radians
 *
 * @param degrees Input in degrees
 * @return Input in radians
 */
public inline f<double> degToRad(double degrees) {
    return degrees * (PI / 180.0);
}

/**
 * Convert radians to degrees
 *
 * @param degrees Input in radians
 * @return Input in degrees
 */
public inline f<double> radToDeg(double radians) {
    return radians * (180.0 / PI);
}

/**
 * Calculate the sine of the input, using the taylor series:
 * sin x = x - x^3/3! + x^5/5! - x^7/7! ...
 *
 * @param x Input number
 * @return Sine of input
 */
public f<double> sin<Numeric>(Numeric x) {
    bool negative = x < 0 ? true : false;
    x = abs(x);
    if x > 360 {
        x -= cast<Numeric>((x / 360) * 360);
    }
    double xRad = degToRad(0.0 + x);
    double res = 0.0;
    double term = 0.0 + xRad;
    double k = 1.0;
    while (res + term != res) {
        res += term;
        k += 2.0;
        term *= -xRad * xRad / k / (k - 1);
    }
    return negative ? -res : res;
}

/**
 * Calculate the cosine of the input, using the taylor series:
 * cos x = 1 - x^2/2! + x^4/4! - x^6/6! ...
 * @param x Input number
 * @return Cosine of input
 */
public f<double> cos<Numeric>(Numeric x) {
    x = abs(x);
    if x > 360 {
        x -= cast<Numeric>((x / 360) * 360);
    }
    double xRad = degToRad(0.0 + x);
    double res = 0.0;
    double term = 1.0;
    double k = 0.0;
    while (res + term != res) {
        res += term;
        k += 2.0;
        term *= -xRad * xRad / k / (k - 1);
    }
    return res;
}

/**
 * Calculate the factorial of the input
 *
 * @param input Input number
 * @return Factorial of input
 */
public inline f<WholeNumber> factorial<WholeNumber>(WholeNumber input) {
    Numeric fac = cast<Numeric>(1);
    for (int i = 1; i <= input; i++) {
        fac *= i;
    }
    return fac;
}
