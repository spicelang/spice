/*ext f<byte*> fopen(string, string);
ext f<int> fclose(byte*);
ext f<int> fputc(int, byte*);
ext f<int> fputs(string, byte*);

f<int> main() {
    byte* file = fopen("./test-file.txt", "w");
    fputs("Hello World!", file);
    fclose(file);
}*/

import "std/io/file";
import "std/type/result";

f<int> main() {
    Result<File> res = openFile("test-file.txt", MODE_WRITE);
    assert res.isOk();
    File file = res.unwrap();
    file.write("test");
    file.close();
}

/*import "../../src-bootstrap/reader/reader";

f<int> main() {
    Reader reader = Reader("./test-file.txt");

    printf("%d", reader.isEOF());
    while !reader.isEOF() {
        printf("%c", reader.getChar());
        reader.advance();
    }
}*/

/*import "std/io/file";

f<int> main() {
    // Write file
    Result<File> fileResult = openFile("./test-file.txt", MODE_WRITE);
    assert fileResult.isOk();
    File file = fileResult.unwrap();
    file.write("Hello, world!\n");
    file.close();

    // Read file
    fileResult = openFile("./test-file.txt", MODE_READ);
    assert fileResult.isOk();
    file = fileResult.unwrap();
    String line = file.readLine();
    printf("%s", line);
    assert line.getRaw() == "Hello, world!\n";
    file.close();

    // Append file
    fileResult = openFile("./test-file.txt", MODE_APPEND);
    assert fileResult.isOk();
    file = fileResult.unwrap();
    file.write("Hello, again!\n");
    file.close();

    // Read file
    fileResult = openFile("./test-file.txt", MODE_READ);
    assert fileResult.isOk();
    file = fileResult.unwrap();
    assert file.readLine() == String("Hello, world!\n");
    assert file.readLine() == String("Hello, again!\n");
    file.close();
}*/