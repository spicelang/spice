#![non.existing.attribute = 22s]