f<bool> isValid(int input = 12) {
    printf("This is a test");
}

f<int> main() {
    bool isValid = isValid();
    printf("Is valid: %d", isValid);
}