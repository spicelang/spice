public type IGlobalResourceManager interface {}