// Imports
import "std/type/int" as intTy;

public type CodeLoc struct {
    unsigned long line
    unsigned long col
    string sourceFilePath
}

public p CodeLoc.ctor(unsigned long line, unsigned long col, string sourceFilePath = "") {
    this.line = line;
    this.col = col;
    this.sourceFilePath = sourceFilePath;
}

/**
 * Returns the code location as a string for using it as a map key or similar
 *
 * @return Code location string
 */
public f<string> toString() {
    return "L" + intTy.toString(line) + "C" + intTy.toString(col);
}

/**
 * Returns the code location in a pretty form
 *
 * @return Pretty code location
 */
public f<string> toPrettyString() {
    if sourceFilePath.empty() {
        return intTy.toString(line) + ":" + intTy.toString(col);
    }
    return sourceFilePath + ":" + intTy.toString(line) + ":" + intTy.toString(col);
}

/**
 * Returns the line number in a pretty form
 *
 * @return Pretty line number
 */
public f<string> toPrettyLine() {
    return "l" + intTy.toString(line);
}