import "std/os/os";
import "std/data/vector";

// Generic types
type T bool|String|int|long|short;

// Enums
type CliOptionMode enum { SET_VALUE, CALL_CALLBACK }

public type CliOption<T> struct {
    string name
    string description
    Vector<string> aliases
    CliOptionMode mode
    T& targetVariable
    p(T&) callback
}

public p CliOption.ctor(string name, T& targetVariable, string description) {
    this.name = name;
    this.description = description;
    this.mode = CliOptionMode::SET_VALUE;
    this.targetVariable = targetVariable;
}

public p CliOption.ctor(string name, p(T&) callback, string description) {
    this.name = name;
    this.description = description;
    this.mode = CliOptionMode::CALL_CALLBACK;
    this.callback = callback;
}

public f<string> CliOption.getName() {
    return this.name;
}

public f<string> CliOption.getDescription() {
    return this.description;
}

public p CliOption.addAlias(string optionName) {
    this.aliases.pushBack(optionName);
}

public f<const Vector<string>&> CliOption.getAliases() {
    return this.aliases;
}

public p CliOption.setTargetValue(T value) {
    if this.mode == CliOptionMode::SET_VALUE {
        this.targetVariable = value;
    }
}

public p CliOption.callCallback(T& value) {
    if this.mode == CliOptionMode::CALL_CALLBACK {
        p(T&) cb = this.callback;
        cb(value);
    }
}