// Link external functions
ext f<string> getenv(string);
ext f<int> putenv(string);

/**
 * Returns the content of an environment variable as string.
 *
 * @return Env variable content or error
 */
public f<Result<string>> getEnv(string name) {
    string value = getenv(name);
    return value != nil<string> ? ok(value) : err<string>(Error("Env var not found"));
}

/**
 * Sets the content of an environment variable to the given value.
 *
 * @return Successful or not
 */
public f<bool> setEnv(string name, string value) {
    String str = String(name);
    str += "=";
    str += value;
    return putenv(str.getRaw()) == 0;
}