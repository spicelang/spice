type T int|dyn|double;

f<int> main() {}