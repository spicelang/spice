import "std/iterators/ranges";

f<int> main() {
    dyn it = range(1, 10);
    assert it.hasNext();
}