type T int|double;

f<T> max<T>(T a, T b) {
    return a > b ? a : b;
}

f<int> main() {
    dyn test = max<short>(1s, 2s);
    printf("Output: %d\n", test);
}