type Driveable interface {
    public p drive(int);
}

type Car struct : Driveable {
    bool driving
}

public p Car.ctor() {
    this.driving = false;
}

public p Car.drive(int param) {
    this.driving = true;
}

f<int> main() {
    Car c = Car();
    Driveable* d = &c;
    d.drive(12);
}

/*import "std/io/cli-parser";

type CliOptions struct {
    bool sayHi = false
}

p callback(bool& value) {
    printf("Callback called with value %d\n", value);
}

f<int> main(int argc, string[] argv) {
    CliParser parser = CliParser("Test Program", "This is a simple test program");
    parser.setVersion("v0.1.0");
    parser.setFooter("Copyright (c) Marc Auberer 2021-2023");

    CliOptions options;
    parser.addFlag("--hi", options.sayHi, "Say hi to the user");
    parser.addFlag("--callback", callback, "Call a callback function");
    parser.addFlag("-cb", p(bool& value) {
        printf("CB called with value %d\n", value);
    }, "Call a callback function");

    parser.parse(argc, argv);

    // Print hi if requested
    if options.sayHi {
        printf("Hi!\n");
    }
}*/

/*type Iterable interface {
    p print();
}

type A struct : Iterable {
    int a
}

p A.print() {
    printf("A: %d\n", this.a);
}

f<int> main() {
    A a = A{5};
    Iterable* i = &a;
    i.print();
}*/