// Std imports
import "std/text/stringstream";

// Ówn imports
import "bootstrap/util/code-loc";

public type ParserErrorType enum {
    PARSING_FAILED,
    NUMBER_OUT_OF_RANGE,
    INVALID_QUALIFIER_COMBINATION,
    INVALID_CHAR_LITERAL,
    INVALID_ATTR_VALUE_TYPE,
    RESERVED_KEYWORD
}

/**
 * Custom exception for errors, occurring while parsing
 */
public type ParserError struct {
    String errorMessage
}

/**
 * Constructor: Used in case that the exact code position where the error occurred is known
 *
 * @param codeLoc Code location where the error occurred
 * @param errorType Type of the error
 * @param message Error message suffix
 */
public p ParserError.ctor(const CodeLoc* codeLoc, const ParserErrorType errorType, const string message) {
    StringStream msg;
    msg << "[Error|Parser] " << codeLoc.toPrettyString() << ": " << this.getMessagePrefix(errorType) << ": " << message;
    this.errorMessage = msg.str();
}

/**
 * Get the prefix of the error message for a particular error
 *
 * @param errorType Type of the error
 * @return Prefix string for the error type
 */
f<string> ParserError.getMessagePrefix(const ParserErrorType errorType) {
    switch errorType {
        case ParserErrorType::PARSING_FAILED: { return "Parsing failed"; }
        case ParserErrorType::NUMBER_OUT_OF_RANGE: { return "Number is out of range"; }
        case ParserErrorType::INVALID_QUALIFIER_COMBINATION: { return "Invalid qualifier combination"; }
        case ParserErrorType::INVALID_CHAR_LITERAL: { return "Invalid char literal"; }
        case ParserErrorType::INVALID_ATTR_VALUE_TYPE: { return "Invalid attribute value type"; }
        case ParserErrorType::RESERVED_KEYWORD: { return "Usage of reserved keyword"; }
        default: { panic(Error("Unknown error")); }
    }
}