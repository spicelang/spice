f<int> main() {
    if 7 {
        printf("Test");
    }
    return 0;
}