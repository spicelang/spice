f<int> main() {
    p(int, int) add = p(int x, int y) {
        return x + y;
    };
}