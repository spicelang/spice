/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/data/vector" as vector;

f<int> main() {
    dyn v = vector.Vector<int>{};
    v.push(4);
    v.push(2);
}*/

//import "os-test2" as s1;
import "std/text/format" as fmt;

f<int> main() {
    /*dyn v1 = s1.Vector<int>{};
    v1.setData<int>(12);
    printf("Data: %d\n", v1.data);

    dyn v2 = s1.Vector<double>{};
    v2.setData<double>(1.5);
    printf("Data: %f\n", v2.data);*/
    printf("%s", fmt.toUpper("test"));
}