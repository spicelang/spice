f<int> main() {
    for int i = 0; i < 15; i++ {
        if i > 6 {
            int j = 6;
            while j > 3 {
                printf("Test");
                break 4;
                j--;
            }
        }
    }
}