f<dyn> testFunction() {
    if true { return "test"; }
    return 0.2;
}

f<int> main() {
    dyn ret = testFunction();
    printf("Result: ", ret);
    return 0;
}