f<int> main() {
    int i;
    i++;
    printf("%d", i);
}