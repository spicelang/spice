import "test1" as test1;

f<int> main() {
    if 1 != 1 {
        printf("If branch");
    } else if 2.0 == 3.1415 {
        printf("Else if 1");
    } else if 2.0 == 2.7183 {
        printf("Else if 2");
    } else {
        printf("Else");
    }
}