import "std/type/int" as i;

f<int> main() {
    bool a = false;
    bool b = true;
    if a = b {
        printf("a: %d, b: %d", a, b);
    } else {
        printf("a: %d, b: %d", a, b);
    }
}

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

/*public f<bool> src(bool x, bool y) {
    return ((x ? 1 : 4) & (y ? 1 : 4)) == 0;
}

public f<int> tgt(int x, int y) {
    return x ^ y;
}

f<int> main() {
    printf("Result: %d, %d", src(false, true), tgt(0, 1));
}*/