const int globalTestVar = 123;