f<int> main() {
    // Plus
    printf("Result: %s\n", String("Hello ") + String("World!"));
    String s1 = String("Hello ");
    printf("Result: %s\n", s1 + " Hi!");
}

/*type Test struct {
    int t
}

p Test.dtor() {
    printf("Dtor called!");
}

f<Test> test() {
    return Test{123};
}

f<int> main() {
   Test t = test();
   printf("%d", t.t);
}*/