type Test struct {
    int f1
    int f2
}

f<int> main() {
    int t = 123;
    switch (t) {
        case 1: {
            printf("1");
        }
        case Test: {
            printf("t");
        }
    }
}