public type IFunction interface {

}
