f<int> main() {
    int i = 123;
    printf("%d", *i);
}