public const int SIZE = 8;
public const byte MIN_VALUE = 0;
public const byte MAX_VALUE = 255;

// Converts a byte to a double
public f<double> toDouble(byte input) {
    return 0.0;
}

// Converts a byte to an int
public f<int> toInt(byte input) {
    return (int) input;
}

// Converts a byte to a short
public f<short> toShort(byte input) {
    return (short) input;
}

// Converts a byte to a long
public f<long> toLong(byte input) {
    return (long) input;
}

// Converts a byte to a char
public f<char> toChar(byte input) {
    return (char) input;
}

// Converts a byte to a string
public f<string> toString(byte input) {
    return "0";
}

// Converts a byte to a bool
public f<bool> toBool(byte input) {
    return input == 1;
}