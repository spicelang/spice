import "std/data/vector";
import "std/data/linked-list";
import "std/math/hash";
import "std/iterator/iterable";
import "std/iterator/iterator";
import "std/data/pair";

// Generic types for key and value
type K dyn;
type V dyn;

type HashEntry<K, V> struct {
    K key
    V value
}

public p HashEntry.ctor(const HashEntry<K, V>& original) {
    this.key = original.key;
    this.value = original.value;
}

public type HashTable<K, V> struct : IIterable<Pair<K, V>> {
    Vector<LinkedList<HashEntry<K, V>>> buckets
}

public p HashTable.ctor(unsigned long bucketCount = 100l) {
    this.buckets = Vector<LinkedList<HashEntry<K, V>>>(bucketCount);
    for unsigned long i = 0l; i < bucketCount; i++ {
        this.buckets.pushBack(LinkedList<HashEntry<K, V>>());
    }
}

/**
 * Insert a key-value pair into the hash table.
 * If the key already exists, the value is updated.
 *
 * @param key The key to insert
 * @param value The value to insert
 */
public p HashTable.upsert(const K& key, const V& value) {
    const LinkedList<HashEntry<K, V>>& bucket = this.getBucket(key);
    foreach const HashEntry<K, V>& entry : bucket {
        if (entry.key == key) {
            entry.value = value;
            return;
        }
    }
    bucket.pushBack(HashEntry<K, V>{key, value});
}

/**
 * Retrieve the value associated with the given key.
 * If the key is not found, panic.
 *
 * @param key The key to look up
 * @return The value associated with the key
 */
public f<V&> HashTable.get(const K& key) {
    foreach const HashEntry<K, V>& entry : this.getBucket(key) {
        if (entry.key == key) {
            return entry.value;
        }
    }
    panic(Error("The provided key was not found"));
}

/**
 * Retrieve the value associated with the given key as Optional<T>.
 * If the key is not found, return an empty optional.
 *
 * @param key The key to look up
 * @return Optional<T>, containing the value associated with the key or empty if the key is not found
 */
public f<Result<V>> HashTable.getSafe(const K& key) {
    foreach const HashEntry<K, V>& entry : this.getBucket(key) {
        if (entry.key == key) {
            return ok(entry.value);
        }
    }
    return err<V>(Error("The provided key was not found"));
}

/**
 * Remove the key-value pair associated with the given key.
 * If the key is not found, do nothing.
 *
 * @param key The key to remove
 */
public p HashTable.remove(const K& key) {
    LinkedList<HashEntry<K, V>>& bucket = this.getBucket(key);
    for unsigned long i = 0l; i < bucket.getSize(); i++ {
        if (bucket.get(i).key == key) {
            bucket.removeAt(i);
            return;
        }
    }
}

/**
 * Check if the hash table contains the given key.
 *
 * @param key The key to check for
 * @return True if the key is found, false otherwise
 */
public f<bool> HashTable.contains(const K& key) {
    foreach const HashEntry<K, V>& entry : this.getBucket(key) {
        if (entry.key == key) {
            return true;
        }
    }
    return false;
}

/**
 * Get the size of the hash table.
 *
 * @return The number of key-value pairs in the hash table
 */
public inline f<unsigned long> HashTable.getSize() {
    result = 0l;
    foreach LinkedList<HashEntry<K, V>>& bucket : this.buckets {
        result += bucket.getSize();
    }
}

/**
 * Checks if the hash table is empty.
 *
 * @return True if empty, false otherwise.
 */
public inline f<bool> HashTable.isEmpty() {
    return this.getSize() == 0l;
}

/**
 * Clear the hash table, removing all key-value pairs.
 */
public inline p HashTable.clear() {
    foreach LinkedList<HashEntry<K, V>>& bucket : this.buckets {
        bucket.clear();
    }
}

inline f<LinkedList<HashEntry<K, V>>&> HashTable.getBucket(const K& key) {
    return this.buckets.get(this.hash(key));
}

inline f<unsigned long> HashTable.hash(const K& key) {
    return hash(key) % this.buckets.getSize();
}

/**
 * Iterator to iterate over a hash table data structure
 */
public type HashTableIterator<K, V> struct : IIterator<Pair<const K&, V&>> {
    HashTable<K, V>& hashTable
    Pair<const K&, V&> currentPair
    unsigned long currentBucketIdx = 0l
    unsigned long currentBucketItemIdx = 0l
    unsigned long cursor = 0l
}

public p HashTableIterator.ctor<K, V>(HashTable<K, V>& hashTable) {
    this.hashTable = hashTable;
    if !this.hashTable.buckets.isEmpty() {
        // Find first bucket that contains any items
        const LinkedList<HashEntry<K, V>>& currentBucket = this.hashTable.buckets.get(this.currentBucketIdx);
        while this.currentBucketIdx + 1 < this.hashTable.buckets.getSize() && currentBucket.isEmpty() {
            currentBucket = this.hashTable.buckets.get(++this.currentBucketIdx);
        }
    }
}

/**
 * Returns the current key-value pair of the hash table
 *
 * @return Current key/value pair
 */
public inline f<Pair<const K&, V&>&> HashTableIterator.get() {
    // Retrieve current bucket
    LinkedList<HashEntry<K, V>>& currentBucket = this.hashTable.buckets.get(this.currentBucketIdx);
    // Retrieve correct entry in the current bucket
    HashEntry<K, V>& hashEntry = currentBucket.get(this.currentBucketItemIdx);
    // Construct pair from key and value
    this.currentPair = Pair<const K&, V&>(hashEntry.key, hashEntry.value);
    return this.currentPair;
}

/**
 * Returns the current index and the current item of the hash table
 *
 * @return Pair of current index and current key/value pair
 */
public inline f<Pair<unsigned long, Pair<const K&, V&>&>> HashTableIterator.getIdx() {
    return Pair<unsigned long, Pair<const K&, V&>&>(this.cursor, this.get());
}

/**
 * Check if the iterator is valid
 *
 * @return true or false
 */
public inline f<bool> HashTableIterator.isValid() {
    // Check if the hash table has no buckets
    if this.hashTable.isEmpty() { return false; }
    // Check if we reached the end of the bucket list
    if this.currentBucketIdx >= this.hashTable.buckets.getSize() { return false; }
    // Check if any more items are to come
    return this.moreItemsAvailable();
}

f<bool> HashTableIterator.moreItemsAvailable() {
    // Are we at the end of the current bucket?
    const LinkedList<HashEntry<K, V>>& currentBucket = this.hashTable.buckets.get(this.currentBucketIdx);
    if this.currentBucketItemIdx + 1 < currentBucket.getSize() {
        return true;
    }
    // Are there more non-empty buckets?
    for unsigned long i = this.currentBucketIdx; i < this.hashTable.buckets.getSize(); i++ {
        const LinkedList<HashEntry<K, V>>& bucket = this.hashTable.buckets.get(i);
        if !bucket.isEmpty() {
            return true;
        }
    }
    return false;
}

p HashTableIterator.moveToNextItem() {
    // Retrieve current bucket
    const LinkedList<HashEntry<K, V>>& currentBucket = this.hashTable.buckets.get(this.currentBucketIdx);
    this.currentBucketItemIdx++;

    // If the current bucket does not contain more items, move to the next bucket that contains items
    if this.currentBucketItemIdx >= currentBucket.getSize() {
        this.currentBucketIdx++;
        if this.currentBucketIdx < this.hashTable.buckets.getSize() {
            currentBucket = this.hashTable.buckets.get(this.currentBucketIdx);
            while this.currentBucketIdx + 1 < this.hashTable.buckets.getSize() && currentBucket.isEmpty() {
                currentBucket = this.hashTable.buckets.get(++this.currentBucketIdx);
            }
        }
        this.currentBucketItemIdx = 0l;
    }
}

/**
 * Moves the cursor to the next key/value pair
 */
public inline p HashTableIterator.next() {
    if !this.isValid() { panic(Error("Calling next() on invalid iterator")); }

    // Move to next item
    this.moveToNextItem();

    // Increment cursor to reflect the current item position
    this.cursor++;
}

/**
 * Retrieve a forward iterator for the hash table
 */
public f<HashTableIterator<K, V>> HashTable.getIterator() {
    return HashTableIterator<K, V>(*this);
}
