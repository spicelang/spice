import "std/io/filepath";
import "std/os/os";

f<int> main() {
    FilePath path = FilePath("C:\Users\Public\Documents");
    path /= "test.txt";
    assert len(path.toString()) == 34;

    printf("All assertions passed!");
}