const int testInt = 0;
double testDouble = 1.5;
string testString = "";
bool testBool = true;
dyn testAuto = false;

4++;

// This is a test comment
f<int> testFunction(double doubleParam) {
    dyn number;
    number = 123;
    result = number | true;

    while testDouble < 2.5 {
        for int i = 12; i < 15; i+=2 {
            return 12;
        }
    }
    return result;
}

p testProcedure(bool boolParam = false, string stringParam) {
    /* Test
    block
    comment */
    double result = testString == "" || testBool ? 5.0 : 1.4;
}