type UnusedInterface interface {
    f<int> testFunction()
}

f<int> main() {}