f<int> main() {
    int testVar = 12;
    {
        printf("Test var: %d\n", testVar);
    }
}