int CONST1 = 123;
int CONST2 = 1234;

f<int> main() {
    printf("1. Constant: %d\n", CONST1);
    printf("2. Constant: %d\n", CONST2);
}