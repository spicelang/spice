// Std imports
import "std/data/vector";
import "std/data/map";

// Own imports
import "bootstrap/ast/ast-nodes";
import "bootstrap/symboltablebuilder/super-type";
import "bootstrap/symboltablebuilder/qual-type";
import "bootstrap/symboltablebuilder/symbol-table-entry";
import "bootstrap/model/generic-type";

// Helper structs
public type Param struct {
    QualType qualType
    bool isOptional = false
}

public type NamedParam struct {
    string name = nil<string>
    QualType qualType
    bool isOptional = false
}

// Type aliases
type ParamList alias Vector<Param>;
type NamedParamList alias Vector<NamedParam>;

public type Function struct {
    String name
    QualType thisType = QualType(SuperType::TY_DYN)
    QualType returnType = QualType(SuperType::TY_DYN)
    ParamList paramList
    Vector<GenericType> templateTypes
    Map<String, QualType> typeMapping
    SymbolTableEntry* entry
    ASTNode* declNode
    bool genericSubstantiation
    bool alreadyTypeChecked
    bool external
    bool used
}