f<int> main() {
    dyn integer = 1;
    printf("%s", &integer);
}