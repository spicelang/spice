f<int> main() {
    double variable;
    printf("Double value: %f", variable);
}