import "std/data/linked-list";

f<int> main() {
    dyn linkedList = LinkedList<int>();
    linkedList.insert(1234);
    linkedList.insert(4567);
    linkedList.insert(7890);
    linkedList.insert(4567);
    linkedList.remove(7890);
}