f<int> main() {
    dyn condition = 1 != 2;
    bool[12] myBoolArray = { condition ? true : false, false, true };

    int i = 2;
    bool itemValue = myBoolArray[i -= 2];
    printf("Value: %u", itemValue);
}