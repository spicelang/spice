type T int|long;

type TestStruct<T> struct {
    T f1
    unsigned long length
}

p TestStruct.ctor(const unsigned long initialLength) {
    length = initialLength;
}

p TestStruct.printLength() {
    printf("%d", this.length);
}

type Alias alias TestStruct<long>;

f<int> main() {
    Alias a = Alias{12345l, 54321l};
    a.printLength();
    dyn b = Alias(12l);
    b.printLength();
}