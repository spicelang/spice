import "std/data/vector";
import "std/data/pair";

f<int> main() {
    Vector<Pair<int, string>> pairVector = Vector<Pair<int, string>>();
    pairVector.pushBack(Pair<int, string>(0, "Hello"));
    pairVector.pushBack(Pair<int, string>(1, "World"));

    Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!\n", p1.getSecond());
}

/*import "std/os/thread";

f<int> fib(int n) {
    if n <= 2 { return 1; }
    return fib(n - 1) + fib(n - 2);
}

p calcFib30() {
    int result = fib(30);
    printf("Thread returned with result: %d\n", result);
}

f<int> main() {
    int threadCount = 8;
    Thread[8] threads = {};
    for unsigned int i = 0; i < threadCount; i++ {
        threads[i] = Thread(calcFib30);
    }
    printf("Started all threads. Waiting for results ...\n");
    for unsigned int i = 0; i < threadCount; i++ {
        Thread& thread = threads[i];
        thread.join();
    }
    printf("Program finished");
}*/

/*type T int|long;

type TestStruct<T> struct {
    T _f1
    unsigned long length
}

p TestStruct.ctor(const unsigned long initialLength) {
    this.length = initialLength;
}

p TestStruct.printLength() {
    printf("%d\n", this.length);
}

type Alias alias TestStruct<long>;

f<int> main() {
    Alias a = Alias{12345l, (unsigned long) 54321l};
    a.printLength();
    dyn b = Alias(12l);
    b.printLength();
}*/

/*type TestStruct struct {
    long lng
    String str
    int i
}

p TestStruct.dtor() {}

f<TestStruct> fct(int& ref) {
    TestStruct ts = TestStruct{ 6l, String("test string"), ref };
    return ts;
}

f<int> main() {
    int test = 987654;
    const TestStruct res = fct(test);
    printf("Long: %d\n", res.lng);
    printf("String: %s\n", res.str.getRaw());
    printf("Int: %d\n", res.i);
}*/