public const int BOOL_SIZE = 1;
public const bool TRUE = true;
public const bool FALSE = false;

// Converts a bool to a double
public f<double> toDouble(bool input) {
    return input ? 1.0 : 0.0;
}

// Converts a bool to an int
public f<int> toInt(bool input) {
    return input ? 1 : 0;
}

// Converts a bool to a short
public f<short> toShort(bool input) {
    return (short) (input ? 1 : 0);
}

// Converts a bool to a long
public f<long> toLong(bool input) {
    return (long) (input ? 1 : 0);
}

// Converts a bool to a byte
public f<byte> toByte(bool input) {
    result = (byte) (input ? 1 : 0);
}

// Converts a bool to a string
public f<string> toString(bool input) {
    return input ? "true" : "false";
}