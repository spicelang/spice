import "std/text/print" as print;
//import "std/runtime/string" as str;

type Test struct {
    int field1
    double field2
}

p Test.ctor() {
    this.field1 = 1;
    this.field2 = 1.0;
}

p Test.dtor() {
    this.field1 = 0;
    this.field2 = 0.0;
}

p Test.setField1(int value) {
    this.field1 = value;
}

f<int> Test.getField1() {
    return this.field1;
}

f<int> main() {
    Test test = Test { 5, 4.567 };
    test.setField1(6);
    print.println("Output:");
    printf("%d", test.getField1());
}