import "source2";

f<int> main() {
    Operand op;
    op++;
}