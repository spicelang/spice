f<int> main() {
    double d;
    len(d);
}