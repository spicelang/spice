// Std imports
import "std/data/vector";
import "std/os/system";

// Own imports
import "../util/memory";

type Base dyn;

public type BlockAllocator<Base> struct {
    IMemoryManager* memoryManager
    Vector<byte*> memoryBlocks
    Vector<Base*> allocatedObjects
    unsigned long blockSize
    unsigned long offsetInBlock = 0l
}

public p BlockAllocator.ctor(IMemoryManager* memoryManager, unsigned long blockSize = 0l) {
    this.memoryManager = memoryManager;
    this.blockSize = blockSize == 0l ? (unsigned long) getPageSize() : blockSize;
    // Allocate the first block
    this.allocateNewBlock();
}

public p BlockAllocator.dtor() {
    // Destruct all objects
    foreach Base* ptr : this.allocatedObjects {
        sDelete(ptr);
    }
    this.allocatedObjects.clear();

    // Free all memory blocks
    foreach byte* block : this.memoryBlocks {
        this.memoryManager.deallocate(block);
    }
    this.memoryBlocks.clear();
}

public p BlockAllocator.allocateNewBlock() {
    // Allocate new block
    heap byte* ptr = this.memoryManager.allocate(this.blockSize);
    if ptr != nil<heap byte*> {
        panic(Error("Could not allocate memory block for BlockAllocator."));
    }

    // Store pointer and reset offset
    this.memoryBlocks.pushBack(ptr);
    this.offsetInBlock = 0l;
}