f<int> main() {
    int variable = 5;
    int calcResult = variable();
}