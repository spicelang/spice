import "std/iterator/iterable";

// Generic type definitions
type T int|long|short;

/**
 * A NumberIterator in Spice can be used to iterate over a range of numbers
 */
public type NumberIterator<T> struct : Iterable<T> {
    T lowerBound // Inclusive
    T upperBound // Inclusive
    unsigned long cursor
}

public p NumberIterator.ctor(T lowerBound, T upperBound) {
    assert lowerBound <= upperBound;
    this.lowerBound = lowerBound;
    this.upperBound = upperBound;
    this.cursor = 0l;
}

/**
 * Check if the number range has another number
 *
 * @return true or false
 */
public inline const f<bool> NumberIterator.hasNext() {
    return this.lowerBound + this.cursor <= this.upperBound;
}

/**
 * Returns the current number of the number range and moves the cursor to the next item
 *
 * @return current item
 */
public inline f<T> NumberIterator.next() {
    assert this.hasNext();
    this.cursor++;
    return (T) (this.lowerBound + this.cursor);
}

/**
 * Returns the current number as well as the current iterator index and moves the cursor
 * to the next item.
 *
 * @return pair of index and item
 */
public inline f<Pair<unsigned long, T>> NumberIterator.nextIdx() {
    assert this.hasNext();
    this.cursor++;
    T currentNumber = (T) (this.lowerBound + this.cursor);
    return Pair<unsigned long, T>(this.cursor, currentNumber);
}

/**
 * Returns the current number of the number range
 */
public inline f<T> NumberIterator.get() {
    return (T) (this.lowerBound + this.cursor);
}

/**
 * Advances the cursor by the given offset
 *
 * @param it NumberIterator
 * @param offset Offset
 */
public inline p operator+=<T>(NumberIterator<T>& it, T offset) {
    it.cursor += offset;
}

/**
 * Move the cursor back by the given offset
 *
 * @param it NumberIterator
 * @param offset Offset
 */
public inline p operator-=<T>(NumberIterator<T>& it, T offset) {
    it.cursor -= offset;
}

/**
 * Convenience wrapper for creating a simple number iterator
 */
public inline f<NumberIterator<T>> range<T>(T begin, T end) {
    return NumberIterator<T>(begin, end);
}