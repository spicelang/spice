p test(int& intRef) {}

f<int> main() {
    test(543210);
}