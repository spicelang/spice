f<int> main() {
    dyn test = "string1" + "string2";
    printf("Test: %s", test);
}