f<int> main() {
    bool b = true;
    foreach string item : b {
        printf("Item: %s", item);
    }
}