type T1 dyn;
type T2 dyn;

inline f<bool> isSame<T1, T2>() {
    return typeid<T1>() == typeid<T2>();
}

f<int> main() {
    assert isSame<int, int>();
    assert !isSame<int, string>();
    assert isSame<double*&, double*&>();
    printf("All assertions passed!\n");
}