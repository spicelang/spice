f<int> main() {
    printf("Test: %d, %f", 3);
}