import "std/iterator/number-iterator";

f<int> main() {
    foreach int i : range(1, 5) {
        printf("%d\n", i);
    }

    /*int[5] testArray = { 1, 6, 3, 11, 5 };
    foreach int idx, int i : array(testArray) {
        printf("%d\n", i);
    }*/


}