import "source1" as s1;

f<int> main() {
    s1::printFormat(1.123);
    s1::printFormat(543);
    s1::printFormat({"Hello", "World"});
}