/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/net/socket" as socket;

f<int> main() {
    socket.Socket s = socket.openServerSocket(8080s, 2);
    printf("Error code: %d", s.errorCode);
    //s.close();
}*/



//import "std/os/threading" as t;
import "std/time/delay" as delay;

f<int> main() {
    printf("Starting one thread ...\n");
    thread -1 {
        delay.delay(500);
        printf("Hello from the thread 1\n");
    }
    thread -1 {
        delay.delay(200);
        printf("Hello from the thread 2\n");
    }
    delay.delay(1000);
    printf("Hello from original\n");
}