// Contains the operating system name in lower case
public const string OS_NAME = "windows";

// Contains the native path separator
public const char PATH_SEPARATOR = '\\';

// System exit codes
public const int EXIT_CODE_SUCCESS = 0;
public const int EXIT_CODE_ERROR = 1;

// Returns true if the current OS is Linux
public f<bool> isLinux() {
    return false;
}

// Returns true  if the current OS is Windows
public f<bool> isWindows() {
    return true;
}

// Returns true  if the current OS is macOS
public f<bool> isMacOS() {
    return false;
}

// Returns true if the current OS is Unix-based
public f<bool> isUnixBased() {
    return false;
}