// File open modes
public const string MODE_READ                 = "r";
public const string MODE_WRITE                = "w";
public const string MODE_APPEND               = "a";
public const string MODE_READ_WRITE           = "r+";
public const string MODE_READ_WRITE_OVERWRITE = "w+";
public const string MODE_READ_WRITE_APPEND    = "a+";
const int O_RDONLY = 0o00000000; // Read only
const int O_WRONLY = 0o00000001; // Write only
const int O_RDWR   = 0o00000002; // Read and write

// Flags for open()
const int O_APPEND    = 0o00002000;  // Set append mode
const int O_ASYNC     = 0o00020000;  // Send a signal when I/O is possible
const int O_CLOEXEC   = 0o02000000;  // Close the file descriptor upon execution of an exec family function
const int O_CREAT     = 0o00000100;  // Create file if it does not exist
const int O_DIRECT    = 0o00040000;  // Prevent file contents from being cached in memory
const int O_DIRECTORY = 0o00200000;  // Fail if not a directory
const int O_DSYNC     = 0o00010000;  // Use synchronized I/O data integrity completion
const int O_EXCL      = 0o00000200;  // Fail if file already exists
const int O_LARGEFILE = 0o00100000;  // Allow large file offsets
const int O_NOATIME   = 0o00020000;  // Do not update file access time
const int O_NOCTTY    = 0o00000400;  // Do not allow control of terminal device
const int O_NOFOLLOW  = 0o00001000;  // Do not follow symlinks
const int O_NONBLOCK  = 0o00004000;  // Use non-blocking I/O
const int O_PATH      = 0o010000000; // Resolve pathname but do not open file
const int O_SYNC      = 0o00004000;  // Use synchronized I/O file integrity completion
const int O_TMPFILE   = 0o020000000; // Create an unnamed temporary file
const int O_TRUNC     = 0o00001000;  // Truncate flag

// File permission modes
public const short S_IRWXU = 0o700s; // Read, write, execute/search by owner
public const short S_IRUSR = 0o400s; // Read permission, owner
public const short S_IWUSR = 0o200s; // Write permission, owner
public const short S_IXUSR = 0o100s; // Execute/search permission, owner
public const short S_IRWXG = 0o070s; // Read, write, execute/search by group
public const short S_IRGRP = 0o040s; // Read permission, group
public const short S_IWGRP = 0o020s; // Write permission, group
public const short S_IXGRP = 0o010s; // Execute/search permission, group
public const short S_IRWXO = 0o007s; // Read, write, execute/search by others
public const short S_IROTH = 0o004s; // Read permission, others
public const short S_IWOTH = 0o002s; // Write permission, others
public const short S_IXOTH = 0o001s; // Execute/search permission, others

// File operation status codes
const int STATUS_OK    = 0;
const int STATUS_ERROR = -1;

// File access flags
const int F_OK = 0; // File existence
const int X_OK = 1; // Can execute
const int W_OK = 2; // Can write
const int R_OK = 4; // Can read

// File seek modes
const int SEEK_SET = 0;
const int SEEK_CUR = 1;
const int SEEK_END = 2;

const int EOF = -1;

type FilePtr alias byte*;

// Link external functions
ext f<FilePtr> fopen(string /*file path*/, string /*mode*/);
ext f<int> fclose(FilePtr /*stream*/);
ext f<int> chmod(string /*file path*/, short /*mode*/);
ext f<int> remove(string /*file path*/);
ext f<int> fgetc(FilePtr /*stream*/);
ext f<int> fputc(int /*char*/, FilePtr /*stream*/);
ext f<int> fputs(string /*string*/, FilePtr /*stream*/);
ext f<int> access(string /*file path*/, int /*mode*/);
ext f<int> fseek(FilePtr /*stream*/, long /*offset*/, int /*whence*/);
ext f<unsigned long> ftell(FilePtr /*stream*/);

public type File struct {
    FilePtr filePtr
    bool isEOF
}

/**
 * Closes the file behind the provided file pointer.
 *
 * @return True if successful, false if not
 */
public f<bool> File.close() {
    result = fclose(this.filePtr) == STATUS_OK;
    this.filePtr = nil<FilePtr>;
}

/**
 * Reads a singe char from the file.
 *
 * @return Char in form of an int, because of EOF = -1.
 */
public f<char> File.readChar() {
    assert !this.isEOF;
    result = (char) fgetc(this.filePtr);
    this.isEOF = result == EOF;
}

/**
 * Reads a single line from the file.
 *
 * @return Line in form of a string
 */
public f<String> File.readLine() {
    assert !this.isEOF;
    result = String();
    char buffer;
    while (buffer = this.readChar()) != EOF {
        if buffer == '\n' { break; }
        result += (char) buffer;
    }
    if buffer == EOF {
        this.isEOF = true;
    }
}

/**
 * Writes a single character to the file.
 *
 * @return True if successful, false if not
 */
public f<bool> File.write(char value) {
    return fputc((int) value, this.filePtr) != STATUS_ERROR;
}

/**
 * Writes a string to the file.
 *
 * @return True if successful, false if not
 */
public f<bool> File.write(string value) {
    return fputs(value, this.filePtr) != STATUS_ERROR;
}

/**
 * Writes a string to the file.
 *
 * @return True if successful, false if not
 */
public f<bool> File.write(String value) {
    return this.write(value.getRaw());
}

/**
 * Returns the size of the file in bytes.
 *
 * @return File size in bytes
 */
public f<unsigned long> File.getSize() {
    // Remember current cursor position
    unsigned long curPos = ftell(this.filePtr);
    // Move the cursor to the end of the file
    fseek(this.filePtr, (long) 0, SEEK_END);
    // Get the cursor position
    unsigned long size = ftell(this.filePtr);
    // Move cursor back to the remembered position
    fseek(this.filePtr, curPos, SEEK_SET);
    return size;
}

/**
 * Checks if the end of the file is reached.
 *
 * @return EOF reached / not reached
 */
public inline f<bool> File.isEOF() {
    return this.isEOF;
}

/**
 * Creates an empty file on disk similar to the 'touch' command on Linux.
 *
 * @return True if successful, false if not
 */
public f<bool> createFile(string path) {
    FilePtr filePtr = fopen(path, MODE_WRITE);
    result = filePtr != nil<FilePtr>;
    fclose(filePtr);
}

/**
 * Changes the permissions of a file.
 *
 * @return True if successful, false if not
 */
public f<bool> changeFilePermissions(string path, short mode) {
    return chmod(path, mode) != STATUS_ERROR;
}

/**
 * Deletes a file from disk.
 *
 * @return True if successful, false if not
 */
public f<bool> deleteFile(string path) {
    return remove(path) == STATUS_OK;
}

/**
 * Opens a (new) file at the specified path with the specified mode.
 *
 * There are predefined constants for the mode available:
 * MODE_READ, MODE_WRITE, MODE_APPEND,
 * MODE_READ_WRITE, MODE_READ_WRITE_OVERWRITE, MODE_READ_WRITE_APPEND
 *
 * @return File pointer
 */
public f<Result<File>> openFile(string path, string mode = MODE_READ) {
    FilePtr fp = fopen(path, mode);
    File file = File{fp, false};
    return fp != nil<FilePtr> ? ok(file) : err<File>(Error("Failed to open file"));
}

/**
 * Reads a whole file from a given path.
 *
 * @return Content in form of a string
 */
public f<Result<String>> readFile(string path) {
    // Open the file in read mode
    Result<File> fileResult = openFile(path, MODE_READ);
    // Check for errors
    if !fileResult.isOk() {
        return err<String>(fileResult.getErr());
    }
    File file = fileResult.unwrap();
    // Read from the file char by char
    char buffer;
    String output = String();
    while (buffer = file.readChar()) != (char) EOF {
        output += (char) buffer;
    }
    // Close the file
    file.close();
    return ok(output);
}

/**
 * Writes a string to a file at a given path.
 *
 * @return True if successful, false if not
 */
public f<Result<bool>> writeFile(string path, string content) {
    // Open the file in write mode
    Result<File> fileResult = openFile(path, MODE_WRITE);
    // Check for errors
    if !fileResult.isOk() {
        return err<bool>(fileResult.getErr());
    }
    File file = fileResult.unwrap();
    // Write the string to the file
    bool success = file.write(content);
    // Close the file
    file.close();
    return ok(success);
}

/**
 * Returns the size of the file at the given paths in bytes.
 *
 * @return File size in bytes
 */
public f<Result<unsigned long>> getFileSize(string path) {
    // Open the file in read mode
    Result<File> fileResult = openFile(path, MODE_READ);
    // Check for errors
    if !fileResult.isOk() {
        return err<unsigned long>(fileResult.getErr());
    }
    File file = fileResult.unwrap();
    // Get the file file
    unsigned long size = file.getSize();
    // Close the file
    file.close();
    return ok(size);
}

/**
 * Checks if a file exists. The function also returns true if the specified path points to a directory.
 *
 * @return Existing / not existing
 */
public f<bool> fileExists(string path) {
    return access(path, F_OK) != STATUS_ERROR;
}

/**
 * Checks if the read permissions to a file are given.
 *
 * @return Readable / not readable
 */
public f<bool> isFileReadable(string path) {
    return access(path, R_OK) != STATUS_ERROR;
}

/**
 * Checks if the write permissions to a file are given.
 *
 * @return Writable / not writable
 */
public f<bool> isFileWritable(string path) {
    return access(path, W_OK) != STATUS_ERROR;
}

/**
 * Checks if the execute permissions to a file are given.
 *
 * @return Executable / not executable
 */
public f<bool> isFileExecutable(string path) {
    return access(path, X_OK) != STATUS_ERROR;
}