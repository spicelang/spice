import "std/data/vector";
import "../../src-bootstrap/bindings/llvm/LLVM" as llvm;

f<int> main() {
    llvm::LLVMContext context;
    llvm::Module module = llvm::Module("test", context);

    llvm::Type returnType;
    Vector<llvm::Type> argTypes;
    llvm::Type funcType = llvm::getFunctionType(returnType, argTypes);
}