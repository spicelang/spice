type T int|long;

type TestStruct<T> struct {
    T f1
    unsigned long length
}

p TestStruct.ctor(const unsigned long initialLength) {
    this.length = initialLength;
}

p TestStruct.printLength() {
    printf("%d\n", this.length);
}

type Alias alias TestStruct<long>;

f<int> main() {
    Alias a = Alias{12345l, 54321l};
    a.printLength();
    dyn b = Alias(12l);
    b.printLength();
}

/*type T string|char;

type TestStruct<T> struct {
    T base
    int test
}

f<int> main() {
    TestStruct<char> s = TestStruct<char>{ 'a', 1 };
    s.printTest();
}

p TestStruct.printTest() {
    printf("Test: %d\n", this.getTest());
}

f<int> TestStruct.getTest() {
    if this.test == 1 {
        this.test++;
        this.printTest();
    }
    return this.test;
}*/

/*ext<byte*> malloc(long);
ext free(byte*);

f<int> main() {
    byte* address = malloc(1l);
    *address = (byte) 12;
    free(address);
}*/

/*f<int> main() {
    int[10] a;
    for int i = 0; i < len(a); i++ {
        a[i] = 1;
    }
    printf("Cell [3]: %d", a[3]);
}*/