f<int> add(int a, int b) {
    return a + b;
}

#[test]
f<bool> testAdd() {
    return false; // Returning false means the test failed
}
