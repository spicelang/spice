// Syscall numbers
public const unsigned short SYSCALL_READ                    = 3us;
public const unsigned short SYSCALL_WRITE                   = 4us;
public const unsigned short SYSCALL_OPEN                    = 5us;
public const unsigned short SYSCALL_CLOSE                   = 6us;
public const unsigned short SYSCALL_WAIT4                   = 7us;
public const unsigned short SYSCALL_LINK                    = 9us;
public const unsigned short SYSCALL_UNLINK                  = 10us;
public const unsigned short SYSCALL_CHDIR                   = 12us;
public const unsigned short SYSCALL_FCHDIR                  = 13us;
public const unsigned short SYSCALL_MKNOD                   = 14us;
public const unsigned short SYSCALL_CHMOD                   = 15us;
public const unsigned short SYSCALL_CHOWN                   = 16us;
public const unsigned short SYSCALL_GETFSSTAT               = 18us;
public const unsigned short SYSCALL_GETDTABLESIZE           = 19us;
public const unsigned short SYSCALL_DUP                     = 20us;
public const unsigned short SYSCALL_PIPE                    = 21us;
public const unsigned short SYSCALL_GETPID                  = 39us;
public const unsigned short SYSCALL_KILL                    = 37us;
public const unsigned short SYSCALL_CREATE                  = 57us;
public const unsigned short SYSCALL_REMOVE                  = 58us;
public const unsigned short SYSCALL_EXECVE                  = 59us;
public const unsigned short SYSCALL_CHDIR_ROOT              = 61us;
public const unsigned short SYSCALL_FCNTL                   = 62us;
public const unsigned short SYSCALL_DUP2                    = 90us;
public const unsigned short SYSCALL_READV                   = 120us;
public const unsigned short SYSCALL_WRITEV                  = 121us;
public const unsigned short SYSCALL_PREAD                   = 140us;
public const unsigned short SYSCALL_PWRITE                  = 141us;
