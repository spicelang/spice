import "std/iterator/number-iterator";

f<int> main() {
    foreach double item : range(1, 5) {
        printf("Item: %f", item);
    }
}