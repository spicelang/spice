import "source3" as s3;

f<int> dummy() {
    return 0;
}