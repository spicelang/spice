// Just a dummy file