import "std/math/fct" as fct;

f<int> main() {
    printf("Abs (int): %d\n", fct::abs(123));
    printf("Abs (int): %d\n", fct::abs(-137));
    printf("Abs (short): %d\n", fct::abs(56s));
    printf("Abs (short): %d\n", fct::abs(-3s));
    printf("Abs (long): %d\n", fct::abs(1234567890l));
    printf("Abs (long): %d\n", fct::abs(-987654321l));
    printf("Abs (double): %f\n", fct::abs(56.123));
    printf("Abs (double): %f\n", fct::abs(-348.12));

    printf("Sin (double): %f\n", fct::sin(78.345));
    printf("Sin (int): %f\n", fct::sin(23));
    printf("Sin (short): %f\n", fct::sin(-68s));
    printf("Sin (long): %f\n", fct::sin(359l));

    printf("Cos (double): %f\n", fct::cos(78.345));
    printf("Cos (int): %f\n", fct::cos(23));
    printf("Cos (short): %f\n", fct::cos(-68s));
    printf("Cos (long): %f\n", fct::cos(359l));
}