// File permission modes
public const int MODE_ALL_RWX   = 0o0000777;
public const int MODE_ALL_RW    = 0o0000666;
public const int MODE_ALL_R     = 0o0000444;

public const int MODE_OWNER_RWX = 0o0000700;
public const int MODE_OWNER_R   = 0o0000400;
public const int MODE_OWNER_W   = 0o0000200;
public const int MODE_OWNER_X   = 0o0000100;

public const int MODE_GROUP_RWX = 0o0000070;
public const int MODE_GROUP_R   = 0o0000040;
public const int MODE_GROUP_W   = 0o0000020;
public const int MODE_GROUP_X   = 0o0000010;

public const int MODE_OTHER_RWX = 0o0000007;
public const int MODE_OTHER_R   = 0o0000004;
public const int MODE_OTHER_W   = 0o0000002;
public const int MODE_OTHER_X   = 0o0000001;

const int F_OK = 0; // File existence
const int X_OK = 1; // Can execute
const int W_OK = 2; // Can write
const int R_OK = 4; // Can read

const int IF_MT          = 61440; // Decimal for octal: 0170000
const int IF_DIR         = 16384; // Decimal for octal: 0040000

const int INVALID_HANDLE = -1; // Decimal for 0xFFFFFFFF

const int FILE_ATTRIBUTE_DIRECTORY = 16;

type FileStat struct {
    unsigned int st_dev    // ID of the device containing file
    unsigned short st_ino  // Inode number
    unsigned short st_mode // File type and mode
    short st_nlink         // Number of hard links
    short st_uid           // User ID of owner
    short st_gid           // Group ID of owner
    unsigned int st_rdev   // Device ID (if special file)
    int st_size            // Total size in bytes
    long st_atime          // Time of last access
    long st_mtime          // Time of last modificatio
    long st_ctime          // Time of last status change
}

type FileTime struct {
    int f1
    int f2
}

type DirEntry struct {
    int fileAttributes
    FileTime f2
    FileTime f3
    FileTime f4
    int f5
    int f6
    int f7
    int f8
    char[260] fileName
    char[14] f9
}

// Link external functions
ext f<int> mkdir(string, int);
ext f<int> rmdir(string);
ext f<int> rename(string, string);
ext f<int> access(string, int);
ext f<int> stat(string, FileStat*);
ext f<byte*> FindFirstFileA(string, DirEntry*) dll;
ext f<bool> FindNextFileA(byte*, DirEntry*) dll;
ext f<bool> FindClose(byte*) dll;

/**
 * Creates an empty directory at the specified path, with the specified mode.
 * Creates at max one directory. If the second last path element does not exist, the operation fails
 *
 * There are predefined constants for the mode available:
 * MODE_ALL_RWX, MODE_ALL_RW, MODE_ALL_R,
 * MODE_OWNER_RWX, MODE_OWNER_R, MODE_OWNER_W, MODE_OWNER_X,
 * MODE_GROUP_RWX, MODE_GROUP_R, MODE_GROUP_W, MODE_GROUP_X,
 * MODE_OTHER_RWX, MODE_OTHER_R, MODE_OTHER_W, MODE_OTHER_X
 *
 * @return Result code of the create operation: 0 = successful, -1 = failed
 */
public f<int> mkDir(string path, int mode) {
    return mkdir(path, mode);
}

/**
 * Creates an empty directory at the specified path, with the specified mode.
 * Unlike mkDir, mkDirs can also create nested path structures.
 *
 * There are predefined constants for the mode available:
 * MODE_ALL_RWX, MODE_ALL_RW, MODE_ALL_R,
 * MODE_OWNER_RWX, MODE_OWNER_R, MODE_OWNER_W, MODE_OWNER_X,
 * MODE_GROUP_RWX, MODE_GROUP_R, MODE_GROUP_W, MODE_GROUP_X,
 * MODE_OTHER_RWX, MODE_OTHER_R, MODE_OTHER_W, MODE_OTHER_X
 *
 * @return Result code of the create operation: 0 = successful, -1 = failed
 */
public f<int> mkDirs(string path, int mode) {
    // ToDo: Implement

    /*char[] pathChars = (char[]) path;
    for int i = 0; i < path.length(); i++ {

    }*/
    return -1;
}

/**
 * Deletes an empty directory at the specified path.
 *
 * @return Result code of the delete operation: 0 = successful, -1 = failed
 */
public f<int> rmDir(string path) {
    return rmdir(path);
}

/**
 * Renames a directory.
 *
 * @return Result code of the rename operation: 0 = successful, -1 = failed
 */
public f<int> renameDir(string oldPath, string newPath) {
    return rename(oldPath, newPath);
}

/**
 * Checks if a directory is existing.
 *
 * @return Existing or not
 */
public f<bool> dirExists(string path) {
    // Check if there exists something, a file or a dir
    if access(path, F_OK) == 0 {
        // Check if it is a dir
        dyn fs = FileStat{};
        if stat(path, &fs) != 0 {
            return false;
        }
        return ((int) fs.st_mode & IF_MT) == IF_DIR;
    }
    return false;
}

/**
 * Lists all files/subdirectories at a given path.
 */
public p listDir(string path) {
    DirEntry dirEntry = DirEntry{};
    byte* handle;
    bool readMore = true;

    // Find first file
    handle = FindFirstFileA(path, &dirEntry);
    if handle == INVALID_HANDLE {
        printf("Dir does not exist\n");
    } else {
        // Read all files
        while readMore {
            printf("Filename: %s\n", dirEntry.fileName);
            // Check if there is another file
            readMore = FindNextFileA(handle, &dirEntry);
        }
    }
    // Close
    FindClose(handle);
}

/**
 * Lists all files/subdirectories at a given path recursively.
 */
public p listDirRecursive(string path) {
    DirEntry dirEntry = DirEntry{};
    byte* handle;
    bool readMore = true;

    // Find first file
    handle = FindFirstFileA(path, &dirEntry);
    if handle == INVALID_HANDLE {
        printf("Dir does not exist\n");
    } else {
        // Read all files
        while readMore {
            printf("Filename: %s\n", dirEntry.fileName);
            if (dirEntry.fileAttributes & FILE_ATTRIBUTE_DIRECTORY) != 0 {
                // ToDo: Uncomment when string concatenation is supported
                //listDirRecursive(path + "\\" + dirEntry.fileName);
            }
            // Check if there is another file
            readMore = FindNextFileA(handle, &dirEntry);
        }
    }
    // Close
    FindClose(handle);
}