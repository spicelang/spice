public f<int> dummy() {
    return 3;
}