import "std/iterator/iterable";
import "std/iterator/iterator";
import "std/data/pair";

type T dyn;

type ExampleContainedType struct {
    int content = 321
}

p ExampleContainedType.ctor(const ExampleContainedType& other) {
    printf("Copy Ctor called!\n");
}

type ExampleIterableType struct : IIterable<ExampleContainedType> {}

type ExampleTypeIterator<T> struct: IIterator<T> {
    T item
    bool isValid = true
}

f<T&> ExampleTypeIterator.get() {
    return this.item;
}

f<Pair<unsigned long, T&>> ExampleTypeIterator.getIdx() {
    return Pair<unsigned long, T&>(0ul, this.item);
}

f<bool> ExampleTypeIterator.isValid() {
    result = this.isValid;
    this.isValid = false;
}

p ExampleTypeIterator.next() {}

f<ExampleTypeIterator<ExampleContainedType>> ExampleIterableType.getIterator() {
    return ExampleTypeIterator<ExampleContainedType>();
}

f<int> main() {
    ExampleIterableType eit;
    foreach ExampleContainedType ct : eit {
        printf("Content: %d\n", ct.content);
    }
}