public type Vector1 struct {
    public int i2
}

public type Vector struct {
    Vector1 i1
}