import "source1";

f<int> main() {
    printf("IsTrue: %d", isTrue());
}