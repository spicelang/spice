// Own imports
import "../lexer/token";

public type Parser struct {

}

public p Parser.ctor(const tk::Token[] tokens, unsigned long tokenCount) {

}

public p Parser.parse() {

}