import "std/iterator/number-iterator";

f<int> main() {
    foreach double i, int item : range(1s, 12s) {
        printf("Item at index %f: %d", i, item);
    }
}