import "std/data/unordered-set";

f<int> main() {
    UnorderedSet<int> unorderedSet;

    // Iterate over empty container
    {
        foreach const int& item : unorderedSet {
            printf("%d\n", item);
        }
    }

    unorderedSet.insert(1);
    unorderedSet.insert(2);
    unorderedSet.insert(3);
    unorderedSet.insert(4);
    unorderedSet.insert(5);
    unorderedSet.insert(99);
    unorderedSet.insert(100);
    unorderedSet.insert(1265);
    unorderedSet.insert(101);
    unorderedSet.insert(102);

    // Iterate over filled container
    foreach const int& item : unorderedSet {
        printf("%d\n", item);
    }
}