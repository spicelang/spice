type Fruit enum {
    BANANA,
    ORANGE
}

f<int> main() {
    printf("Test: %d", Fruit::ORANGE);
}