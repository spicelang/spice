f<int> main() {
    f<string>() callbackWithoutArgs = f<string>() {
        return "Callback called!\n";
    };
    printf("%s", callbackWithoutArgs());

    f<bool>(String&, double) callbackWithArgs1 = f<bool>(String& str, double d) {
        printf("Callback called with args: %s, %f\n", str, d);
        return str.getRaw() == "Hello" && d == 3.14;
    };
    printf("%d\n", callbackWithArgs1(String("Hello"), 3.14));

    f<short>(String, short) callbackWithArgs2 = f<short>(String str, short b) {
        printf("Callback called with args: %s, %d\n", str, b);
        return ~b;
    };
    printf("%d\n", (callbackWithArgs2(String("Hello World!"), 321s) ^ 956s) == 1 ? 9 : 12);
}

/*f<int> main() {
    int z = 2;
    int w = 3;
    p(int&) foo = p(int& x) { // {ptr (fctPtr), ptr (captureStructPtr)}
        //x += z + w;
        x = 5;
    };
    int x = 1;
    foo(x); // Load fctPtr and call it with captureStructPtr
    printf("%d", x);
}*/

/*type T int|long;

type TestStruct<T> struct {
    T _f1
    unsigned long length
}

p TestStruct.ctor(const unsigned long initialLength) {
    this.length = initialLength;
}

p TestStruct.printLength() {
    printf("%d\n", this.length);
}

type Alias alias TestStruct<long>;

f<int> main() {
    Alias a = Alias{12345l, (unsigned long) 54321l};
    a.printLength();
    dyn b = Alias(12l);
    b.printLength();
}*/

/*type TestStruct struct {
    long lng
    String str
    int i
}

p TestStruct.dtor() {}

f<TestStruct> fct(int& ref) {
    TestStruct ts = TestStruct{ 6l, String("test string"), ref };
    return ts;
}

f<int> main() {
    int test = 987654;
    const TestStruct res = fct(test);
    printf("Long: %d\n", res.lng);
    printf("String: %s\n", res.str.getRaw());
    printf("Int: %d\n", res.i);
}*/