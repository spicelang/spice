public const unsigned int DOUBLE_SIZE = 64;
public const double DOUBLE_MIN_VALUE = -1.7976931348623157e+308;
public const double DOUBLE_MAX_VALUE = 1.7976931348623157e+308;

ext f<unsigned int> snprintf(char*, unsigned long, string, double);

// Converts a double to an int
public f<int> toInt(double input) {
    return cast<int>(input);
}

// Converts a double to a short
public f<short> toShort(double input) {
    return cast<short>(input);
}

// Converts a double to a long
public f<long> toLong(double input) {
    return cast<long>(input);
}

// Converts a double to a string
public f<String> toString(double input) {
    const unsigned int length = snprintf(nil<char*>, 0l, "%f", input);
    result = String(length); // Assuming this length is enough
    snprintf(cast<char*>(result.getRaw()), length + 1l, "%f", input);
}

// Converts a double to a boolean
public f<bool> toBool(double input) {
    return input >= 0.5;
}