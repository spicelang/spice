f<bool> condFct() {
    return false;
}

f<string> trueFct() {
    assert false; // Should not be called
    return "true";
}

f<string> falseFct() {
    return "false";
}

f<int> main() {
    printf("Result: %s", condFct() ? trueFct() : falseFct());
}