type Nested struct {
    string nested1
    bool* nested2
}

type TestStruct struct {
    signed int* field1
    double field2
    Nested* nested
}

f<int> main() {
    int input = 12;
    bool boolean = true;
    Nested nestedInstance = Nested { "Hello World!", &boolean };
    dyn instance = TestStruct { &input, 46.34, &nestedInstance };
    TestStruct instance1 = instance;
    printf("Field1: %d, field2: %f", *instance.nested.nested2, instance1.field2);
    printf("Output: %s, %p", instance1.nested.nested1, instance.field1);
}