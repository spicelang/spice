type T int|double|short|long;
type U bool[]|int[];

f<int> sumNumbers<T>(T[] numberArray, long arrayLength) {
    result = 0;
    for long i = 0l; i < arrayLength; i++ {
        result += numberArray[i];
    }
}

p printData<U>(long arrayLength, U list) {
    for long i = 0l; i < arrayLength; i++ {
        printf("Data: %d\n", list[i]);
    }
}

f<int> main() {
    short[7] numberList1 = [ 1s, 2s, 3s, 4s, 5s, 6s, 7s ];
    int result1 = sumNumbers(numberList1, len(numberList1));

    long[4] numberList2 = [ 10l, 12l, 14l, 16l ];
    int result2 = sumNumbers(numberList2, len(numberList2));

    dyn resultList = [result1, result2];
    printData(len(resultList), resultList);

    printf("Results: %d, %d\n", result1, result2);
}