// Imports
import "std/text/print";
import "std/data/pair";
import "./driver";
import "./global/global-resource-manager";
import "./ast/ast-nodes";

type CompileStageType enum {
    NONE,
    LEXER,
    PARSER,
    CST_VISUALIZER,
    AST_BUILDER,
    AST_OPTIMIZER,
    AST_VISUALIZER,
    IMPORT_COLLECTOR,
    SYMBOL_TABLE_BUILDER,
    TYPE_CHECKER_PRE,
    TYPE_CHECKER_POST,
    IR_GENERATOR,
    IR_OPTIMIZER,
    OBJECT_EMITTER
}

type CompileStageIOType enum {
    IO_CODE,
    IO_TOKENS,
    IO_CST,
    IO_AST,
    IO_IR,
    IO_OBJECT_FILE
}

type TimerOutput struct {
  unsigned long lexer = 0l
  unsigned long parser = 0l
  unsigned long cstVisualizer = 0l
  unsigned long astBuilder = 0l
  unsigned long astVisualizer = 0l
  unsigned long importCollector = 0l
  unsigned long symbolTableBuilder = 0l
  unsigned long typeCheckerPre = 0l
  unsigned long typeCheckerPost = 0l
  unsigned long irGenerator = 0l
  unsigned long irOptimizer = 0l
  unsigned long objectEmitter = 0l
  unsigned long executionEngine = 0l
}

/**
 * Collects the output of the compiler for debugging
 */
type CompilerOutput struct {
    String cstString
    String astString
    String symbolTableString
    String irString
    String irOptString
    String asmString
    Vector<CompilerWarning> warnings
    TimerOutput times
}

type NameRegistryEntry struct {
    String name
    SymbolTableEntry* targetEntry
    Scope* targetScope
    SymbolTableEntry* importEntry
    String predecessorName
}

/**
 * Represents a single source file
 */
public type SourceFile struct {
    public String name
    public String fileName
    public String filePath
    public String fileDir
    public String objectFilePath
    public bool stdFile = false
    public bool mainFile = true
    public CompilerOutput compilerOutput
    public SourceFile* parent
    public String cacheKey
    public bool restoredFromCache = false
    public EntryNode ast
    public Scope globalScope
    //public llvm::Module llvmModule
    public Map<String, Pair<SourceFile, const ASTNode*>> dependencies
    public Map<String, NameRegistryEntry> exportedNameRegistry

    GlobalResourceManager& resourceManager
    unsigned short importedRuntimeModules = 0s
    unsigned short totalTypeCheckerRuns = 0s
}

public p SourceFile.ctor(GlobalResourceManager &resourceManager, SourceFile* parent, const String& name, const String& filePath, bool stdFile) {
    // Copy data
    this.resourceManager = resourceManager;
    this.parent = parent;
    this.name = name;
    this.filePath = filePath;
    this.stdFile = stdFile;

    // Deduce fileName and fileDir
    /*this.fileName = ;
    this.fileDir = ;*/
}

public p SourceFile.runLexer() {
    // Lex this source file
}

public p SourceFile.runParser() {
    // Parse this source file
}

public p SourceFile.runCSTVisualizer(string* output) {
    // Only execute if enabled
    if !cliOptions.dumpCST && !cliOptions.testMode { return; }

    // ToDo: Extend
}

public p SourceFile.runASTBuilder() {
    // Transform the imported source files
    // ToDo: Extend
}

public p SourceFile.runASTVisualizer(string* output) {
    // Only execute if enabled
    if !cliOptions.dumpAST && !cliOptions.testMode { return; }

    // ToDo: Extend
}

public p SourceFile.runImportCollector() {

}

public p SourceFile.runSymbolTableBuilder() {

}

public p SourceFile.runTypeChecker() {

}

p SourceFile.runTypeCheckerPre() {

}

p SourceFile.runTypeCheckerPost() {

}

public p SourceFile.runIRGenerator() {

}

public p SourceFile.runDefaultIROptimizer() {

}

public p SourceFile.runObjectEmitter() {

}

public p SourceFile.concludeCompilation() {

}

public p SourceFile.runFrontEnd() {

}

public p SourceFile.runMiddleEnd() {

}

public p SourceFile.runBackEnd() {

}

f<bool> SourceFile.isAlreadyImported(const String& filePathSearch) {
    // Check if the current source file corresponds to the path to search
    if this.filePath == filePathSearch { return true; }
    // Check parent recursively
    return this.parent != nil<SourceFile*> && this.parent.isAlreadyImported(filePathSearch);
}