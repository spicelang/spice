f<int> main() {
    dyn var;
    printf("Test %d", var);
}