import "std/text/format";

f<int> main() {
    printf("toUpper: %c\n", toUpper('j'));
    printf("toUpper: %s\n", toUpper(String("This is a test.")));
    printf("toLower: %c\n", toLower('L'));
    printf("toLower: %s\n", toLower(String("This is a test.")));
    printf("capizalize: %s\n", capitalize(String("word")));

    printf("formatStorageSize: %s\n", formatStorageSize(1l));
    printf("formatStorageSize: %s\n", formatStorageSize(1l, true));
    printf("formatStorageSize: %s\n", formatStorageSize(1234l));
    printf("formatStorageSize: %s\n", formatStorageSize(1234l, true));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567l));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567l, true));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567890l));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567890l, true));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567890123l));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567890123l, true));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567890123456l));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567890123456l, true));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567890123456789l));
    printf("formatStorageSize: %s\n", formatStorageSize(1234567890123456789l, true));
}