f<dyn> calledFunction(int mandatoryParam, dyn optionalParam = true) {
    printf("Mandatory: %d", mandatoryParam);
    printf("Optional: %d", optionalParam);
    return 0.1;
}

f<int> main() {
    dyn res = calledFunction(1, false);
    printf("Result: %d", res);
    return 0;
}