// Constants
const unsigned long INITIAL_ALLOC_COUNT = 5l;
const unsigned int RESIZE_FACTOR = 2;

// Link external functions
ext<byte*> malloc(long);
ext<byte*> realloc(byte*, int);
ext free(byte*);
ext<byte*> memcpy(byte*, byte*, int);

// Add generic type definition
type T dyn;

/**
 * A stack in Spice is a commonly used data structure, which uses the FiLo (first in, last out) principle.
 *
 * Time complexity:
 * Insert: O(1)
 * Delete: O(1)
 * Search: O(n)
 *
 * Stacks pre-allocate space using an initial size and a resize factor to not have to re-allocate
 * with every item pushed.
 */
public type Stack<T> struct {
    T* contents             // Pointer to the first data element
    unsigned long capacity  // Allocated number of items
    unsigned long size      // Current number of items
}

public p Stack.ctor(unsigned long initAllocItems, const T &defaultValue) {
    // Allocate space for the initial number of elements
    this.ctor(initAllocItems);
    // Fill in the default values
    for unsigned long index = 0; index < initAllocItems; index++ {
        unsafe {
            this.contents[index] = defaultValue;
        }
    }
    this.size = initAllocItems;
}

public p Stack.ctor(unsigned int initAllocItems) {
    this.ctor((unsigned long) initAllocItems);
}

public p Stack.ctor(unsigned long initAllocItems = INITIAL_ALLOC_COUNT) {
    // Allocate space for the initial number of elements
    const long itemSize = sizeof(type T) / 8l;
    unsafe {
        this.contents = (T*) malloc(itemSize * initAllocItems);
    }
    this.size = 0l;
    this.capacity = initAllocItems;
}

public p Stack.dtor() {
    // Free all the memory
    unsafe {
        free((byte*) this.contents);
    }
}

/**
 * Add an item to the stack
 */
public p Stack.push(const T& item) {
    // Check if we need to re-allocate memory
    if this.isFull() {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Insert the element at the back
    unsafe {
        this.contents[(int) this.size++] = item;
    }
}

/**
 * Retrieve item and remove it from the stack
 */
public f<T&> Stack.pop() {
    // Pop the element from the stack
    unsafe {
        return this.contents[(int) --this.size];
    }
}

/**
 * Retrieve the current size of the stack
 *
 * @return Current size of the stack
 */
public f<long> Stack.getSize() {
    return this.size;
}

/**
 * Retrieve the current capacity of the stack
 *
 * @return Current capacity of the stack
 */
 public f<long> Stack.getCapacity() {
     return this.capacity;
 }

/**
 * Checks if the queue contains any items at the moment
 *
 * @return Empty or not empty
 */
public f<bool> Stack.isEmpty() {
    return this.size == 0;
}

/**
 * Checks if the queue exhausts its capacity and needs to resize at the next call of push
 *
 * @return Full or not full
 */
public f<bool> Stack.isFull() {
    return this.size == this.capacity;
}

/**
 * Frees allocated memory that is not used by the queue
 */
public p Stack.pack() {
    // Return if no packing is required
    if this.isFull() { return; }
    // Pack the array
    this.resize(this.size);
}

/**
 * Re-allocates heap space for the queue contents
 */
p Stack.resize(unsigned long itemCount) {
    // Allocate the new memory
    const long itemSize = sizeof(type T) / 8l;
    unsafe {
        byte* oldAddress = (byte*) this.contents;
        int newSize = (int) (itemSize * itemCount);
        T* newMemory = (T*) realloc(oldAddress, newSize);
        this.contents = newMemory;
    }
    // Set new capacity
    this.capacity = itemCount;
}