// Imports
import "Token" as tk;