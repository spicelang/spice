f<int> main() {
    return 0;
}

f<int> main() {
    return 1;
}