// Std imports
import "std/type/any";

public type IAbstractAstVisitor interface {
    f<Any> visitEntry(EntryNode*);
    f<Any> visitMainFctDef(EntryNode*);
    f<Any> visitFctDef(EntryNode*);
    f<Any> visitProcDef(EntryNode*);
}