//import "std/os/os" as os;

// File permission modes
const int MODE_ALL_RWX   = 511;   // Decimal for octal: 0000777
const int MODE_ALL_RW    = 438;   // Decimal for octal: 0000666
const int MODE_ALL_R     = 292;   // Decimal for octal: 0000444

const int MODE_OWNER_RWX = 448;   // Decimal for octal: 0000700
const int MODE_OWNER_R   = 256;   // Decimal for octal: 0000400
const int MODE_OWNER_W   = 128;   // Decimal for octal: 0000200
const int MODE_OWNER_X   = 64;    // Decimal for octal: 0000100

const int MODE_GROUP_RWX = 56;    // Decimal for octal: 0000070
const int MODE_GROUP_R   = 32;    // Decimal for octal: 0000040
const int MODE_GROUP_W   = 16;    // Decimal for octal: 0000020
const int MODE_GROUP_X   = 8;     // Decimal for octal: 0000010

const int MODE_OTHER_RWX = 7;     // Decimal for octal: 0000007
const int MODE_OTHER_R   = 4;     // Decimal for octal: 0000004
const int MODE_OTHER_W   = 2;     // Decimal for octal: 0000002
const int MODE_OTHER_X   = 1;     // Decimal for octal: 0000001

const int F_OK = 0; // File existence
const int X_OK = 1; // Can execute
const int W_OK = 2; // Can write
const int R_OK = 4; // Can read

const int IF_DIR         = 16384; // Decimal for octal: 0040000

type FileStat struct {
    int f1
    short f2
    short st_mode
    short f4
    short f5
    short f6
    int f7
    int f8
    long f9
    long f10
    long f11
}

// Link external functions
ext<int> mkdir(char*, int);
ext<int> rmdir(char*);
ext<int> rename(char*, char*);
ext<int> access(char*, int);
ext<int> stat(char*, FileStat*);

/**
 * Creates an empty directory at the specified path, with the specified mode.
 * Creates at max one directory. If the second last path element does not exist, the operation fails
 *
 * There are predefined constants for the mode available:
 * MODE_ALL_RWX, MODE_ALL_RW, MODE_ALL_R,
 * MODE_OWNER_RWX, MODE_OWNER_R, MODE_OWNER_W, MODE_OWNER_X,
 * MODE_GROUP_RWX, MODE_GROUP_R, MODE_GROUP_W, MODE_GROUP_X,
 * MODE_OTHER_RWX, MODE_OTHER_R, MODE_OTHER_W, MODE_OTHER_X
 *
 * @return Result code of the create operation: 0 = successful, -1 = failed
 */
f<int> mkDir(string path, int mode) {
    return mkdir((char*) path, mode);
}

/**
 * Creates an empty directory at the specified path, with the specified mode.
 * Unlike mkDir, mkDirs can also create nested path structures.
 *
 * There are predefined constants for the mode available:
 * MODE_ALL_RWX, MODE_ALL_RW, MODE_ALL_R,
 * MODE_OWNER_RWX, MODE_OWNER_R, MODE_OWNER_W, MODE_OWNER_X,
 * MODE_GROUP_RWX, MODE_GROUP_R, MODE_GROUP_W, MODE_GROUP_X,
 * MODE_OTHER_RWX, MODE_OTHER_R, MODE_OTHER_W, MODE_OTHER_X
 *
 * @return Result code of the create operation: 0 = successful, -1 = failed
 */
f<int> mkDirs(string path, int mode) {
    // ToDo: Implement

    /*char[] pathChars = (char[]) path;
    for int i = 0; i < path.length(); i++ {

    }*/
    return -1;
}

/**
 * Deletes an empty directory at the specified path.
 *
 * @return Result code of the delete operation: 0 = successful, -1 = failed
 */
f<int> rmDir(string path) {
    return rmdir((char*) path);
}

/**
 * Renames a directory.
 *
 * @return Result code of the rename operation: 0 = successful, -1 = failed
 */
f<int> renameDir(string oldPath, string newPath) {
    return rename((char*) oldPath, (char*) newPath);
}

/**
 * Checks if a directory is existing.
 *
 * @return Existing or not
 */
f<bool> dirExists(string path) {
    printf("Testing ...");
    // Check if there exists something, a file or a dir
    int accessResult = access((char*) path, F_OK);
    printf("Access result: %d", accessResult);
    if accessResult == 0 {
        prinf("Found something")
        // Check if it is a dir
        dyn fs = new FileStat {};
        stat((char*) path, &fs);
        prinf("Test: %d\n", fs.st_mode)
        return ((int) fs.st_mode & IF_DIR) == 1;
    }
    prinf("Not found at all")
    return false;
}