p testProc(int[]** nums) {
    int[] nums1 = **nums;
    nums1[2] = 10;
    printf("1: %d\n", nums1[0]);
    printf("2: %d\n", nums1[1]);
    printf("3: %d\n", nums1[2]);
    printf("4: %d\n", nums1[3]);
}

f<int> main() {
    int[4] intArray = { 1, 2, 3, 4 };
    printf("1: %d\n", intArray[1]);
    testProc(& &intArray);

    string test = "test";
    char c1 = test[2];
    printf("Char: %c\n", c1);
}