import "../../src-bootstrap/lexer/Reader.spice";

f<int> main() {
    Reader reader = Reader("./test.spice");

}