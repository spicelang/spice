type TestStruct struct {
    int field1
    double field2
}

f<int> main() {
    int input = 12;
    TestStruct instance = new TestStruct { input, 46.34 };
    //printf("Field1: %d, field2: %f", instance.field1, instance.field2);
}