f<int> main() {
    String s = String("Hello ");
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.append("World!");
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.append('?');
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.append('!');
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    printf("Equals: %d\n", s.opEquals("Hello World!?!"));
    printf("Equals: %d\n", s.opEquals("Hello World!!"));
    printf("Not Equals: %d\n", s.opNotEquals("Hello World!?!"));
    printf("Not Equals: %d\n", s.opNotEquals("Hello World!!"));
    s.clear();
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s.reserve(100l);
    printf("Content: %s\n", s.getRaw());
    printf("Length: %d\n", s.getLength());
    printf("Capacity: %d\n\n", s.getCapacity());
    s = String("");
    printf("Empty: %d\n", s.isEmpty());
    s.append('a');
    printf("Empty: %d", s.isEmpty());
}