/**
 * Check if a short is a power of two
 *
 * @param input Input number
 * @return Is power of two
 */
public f<bool> isPowerOfTwo(short input) {
    return (input & (input - 1s)) == 0s;
}