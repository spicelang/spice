f<int> main() {
    int test = "Test";
    return 0;
}