import "../../src-bootstrap/parser/parser";

f<int> main() {
    Lexer lexer = Lexer("./text-file.spice");
    Parser parser = Parser(lexer);
    parser.parse();
}