/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/net/socket" as socket;

f<int> main() {
    socket.Socket s = socket.openServerSocket(8080s, 2);
    printf("Error code: %d", s.errorCode);
    //s.close();
}*/

f<int> fib(int n) {
    if n <= 2 { return 1; }
    return fib(n - 1) + fib(n - 2);
}

f<int> main() {
    int threadCount = 8;
    byte*[8] threads = {};
    for int i = 0; i < threadCount; i++ {
        threads[i] = thread {
            int result = fib(46);
            printf("Thread %d returned with result: %d\n", tid(), result);
        };
    }
    printf("Started all threads. Waiting for results ...\n");

    join(threads);

    printf("Program finished");
}