import "bootstrap/bindings/llvm/llvm" as llvm;
import "std/data/vector";

f<int> main() {
    llvm::initializeNativeTarget();
    llvm::initializeNativeAsmPrinter();

    heap string targetTriple = llvm::getDefaultTargetTriple();
    string error;
    llvm::Target target = llvm::getTargetFromTriple(targetTriple, &error);
    llvm::TargetMachine targetMachine = target.createTargetMachine(targetTriple, "generic", "", llvm::LLVMCodeGenOptLevel::Default, llvm::LLVMRelocMode::Default, llvm::LLVMCodeModel::Default);

    llvm::LLVMContext context;
    llvm::Module module = llvm::Module("test", context);
    module.setDataLayout(targetMachine.createDataLayout());
    //module.setTargetTriple(targetTriple); // This emits target dependent information in the IR, which is not what we want here.
    llvm::Builder builder = llvm::Builder(context);

    llvm::Type returnType = builder.getInt32Ty();
    Vector<llvm::Type> argTypes;
    llvm::Type funcType = llvm::getFunctionType(returnType, argTypes);
    llvm::Function func = llvm::Function(module, "main", funcType);
    func.setLinkage(llvm::LLVMLinkage::ExternalLinkage);

    llvm::BasicBlock entry = llvm::BasicBlock(context, "");
    func.pushBack(entry);
    builder.setInsertPoint(entry);

    llvm::Value calcResult = builder.createAdd(builder.getInt32(1), builder.getInt32(2), "calcResult");

    llvm::Value helloWorldStr = builder.createGlobalStringPtr("Hello, world!\n", "helloWorldStr");
    Vector<llvm::Type> printfArgTypes;
    printfArgTypes.pushBack(builder.getPtrTy());
    printfArgTypes.pushBack(builder.getInt32Ty());
    llvm::Type printfFuncType = llvm::getFunctionType(builder.getInt32Ty(), printfArgTypes, true);
    llvm::Function printfFunc = module.getOrInsertFunction("printf", printfFuncType);

    Vector<llvm::Value> printfArgs;
    printfArgs.pushBack(helloWorldStr);
    printfArgs.pushBack(calcResult);
    builder.createCall(printfFunc, printfArgs);

    builder.createRet(builder.getInt32(0));

    assert !llvm::verifyFunction(func);
    string output;
    assert !llvm::verifyModule(module, &output);

    printf("%s", module.print());
}