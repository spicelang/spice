// Constants
const unsigned long INITIAL_ALLOC_COUNT = 5l;
const unsigned int RESIZE_FACTOR = 2;

// Link external functions
ext f<byte*> malloc(long);
ext f<byte*> realloc(byte*, int);
ext p free(byte*);
ext f<byte*> memcpy(byte*, byte*, int);

// Add generic type definitions
type K dyn;
type V dyn;

/**
 * A map in Spice is a commonly used data structure, which can be used to represent a list of key value pairs.
 *
 * Time complexity:
 * Insert: O(1)
 * Delete:
 * Search: O(1)
 */
public type Map<K, V> struct {

}

public p Map.ctor() {

}