f<int> main() {
    // Directly
    printf("%d\n", String("").isEmpty());
    printf("%d\n", String("Hello").isEmpty());
    printf("%d\n", String("Hello!").getLength());
    printf("%d\n", String("Hello World!").getLength());
    printf("%d\n", String("Hello!").getCapacity());
    printf("%d\n", String("Hello World!").getCapacity());
    printf("%d\n", String("Hello").isFull());
    printf("%d\n", String("Hello World!").isFull());
    printf("%d\n", String("Hello World!").find("ell"));
    printf("%d\n", String("Hello World!").find("Wort"));
    printf("%d\n", String("Hello World!").find("H"));
    printf("%d\n", String("Hello World!").find("!"));
    printf("%d\n", String("Hello World!").find(" ", 12));
    printf("%d\n", String("Hello World!").contains("abc"));
    printf("%d\n", String("Hello World!").contains("Hello"));
    printf("%d\n", String("Hello World!").contains("World!"));
    printf("%d\n", String("Hello World!").contains("o W"));
}

/*f<int> main() {
    String testString;
    printf("Test: %s\n", testString);
    testString += "Hi!";
    printf("Test: %s\n", testString);
    //testString = String("Lorem ipsum dolor sit amet, consetetur sadipscing elitr, sed diam nonumy eirmod tempor invidunt ut labore et dolore magna aliquyam erat, sed diam voluptua. At vero eos et accusam et justo duo dolores et ea rebum. Stet clita kasd gubergren, no sea takimata sanctus est Lorem ipsum dolor sit amet. Lorem ipsum dolor sit amet, consetetur sadipscing elitr, sed diam nonumy eirmod tempor invidunt ut labore et dolore magna aliquyam erat, sed diam voluptua. At vero eos et accusam et justo duo dolores et ea rebum. Stet clita kasd gubergren, no sea takimata sanctus est Lorem ipsum dolor sit amet.");

    //printf("Length: %d\n", testString.getLength());
    //printf("Capacity: %d", testString.getCapacity());
}*/

/*f<int> main() {
    String s = String("Hello ");
    printf("Output: %s\n", s);
    s = String("");
    printf("Output: %s\n", s);
}*/

/*type Visitor struct {

}

type SymbolTable struct {

}

type VisitableNode interface {
    f<bool> accept(Visitor*)
}

type AstNode struct : VisitableNode {

}

f<bool> AstNode.accept(Visitor* v) {
    return true;
}

type AstEntryNode struct : VisitableNode {
    AstNode astNode
    SymbolTable* fctScope
    bool hasArgs
}

f<bool> AstEntryNode.accept(Visitor* v) {
    return true;
}

f<int> main() {
    dyn entryNode = AstEntryNode{};
    printf("%d", entryNode.hasArgs);
}*/

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

/*public f<bool> src(bool x, bool y) {
    return ((x ? 1 : 4) & (y ? 1 : 4)) == 0;
}

public f<int> tgt(int x, int y) {
    return x ^ y;
}

f<int> main() {
    printf("Result: %d, %d", src(false, true), tgt(0, 1));
}*/