f<int> main() {
    // Directly
    printf("%d\n", "".isEmpty());
    printf("%d\n", "Hello".isEmpty());
    printf("%d\n", "Hello!".getLength());
    printf("%d\n", "Hello World!".getLength());
    printf("%d\n", "Hello!".getCapacity());
    printf("%d\n", "Hello World!".getCapacity());
    printf("%d\n", "Hello".isFull());
    printf("%d\n", "Hello World!".isFull());

    // Via variable
    string var = "";
    printf("%d\n", var.isEmpty());
    var = "Hello";
    printf("%d\n", var.isEmpty());
    var = "Hello!";
    printf("%d\n", var.getLength());
    var = "Hello World!";
    printf("%d\n", var.getLength());
    var = "Hello!";
    printf("%d\n", var.getCapacity());
    var = "Hello World!";
    printf("%d\n", var.getCapacity());
}