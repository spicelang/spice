type Person struct {
    string* firstName
    string* lastName
    int age
}

type Person struct {
    int age
    double* height
}

f<int> main() {}