type Person interface {
    f<int> dump();
}

type Person interface {
    p print();
}

f<int> main() {}