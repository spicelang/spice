// See Issue #155 (fixed)

type T dyn;

public type Vector<T> struct {
    T* contents
    unsigned long capacity
    unsigned long size
    unsigned int itemSize
}

public f<int> Vector.get(long index) {
    if (index <= size) { // size instead this.size
        return 1;
    }
    return 0;
}

f<int> main() {
    dyn v = Vector<int>{};
    int v0 = v.get(0l);
}

/*import "std/net/http" as http;

f<int> main() {
    http::HttpServer server = http::HttpServer();
    server.serve("/test", "Hello World!");
}*/

/*public f<bool> src(bool x, bool y) {
    return ((x ? 1 : 4) & (y ? 1 : 4)) == 0;
}

public f<int> tgt(int x, int y) {
    return x ^ y;
}

f<int> main() {
    printf("Result: %d, %d", src(false, true), tgt(0, 1));
}*/