f<int> add(int a, int b) {
    return a + b;
}

#[test=true, test.name="Test for add function", test.skip=false]
f<bool> testAdd() {
    assert add(1, 2) == 3;
    assert add(2, 2) == 4;
    assert add(3, 2) == 5;

    return true;
}

f<int> main() {
    printf("%d\n", add(1, 2));
}
