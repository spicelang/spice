/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec.Vector<pair.Pair<int, string>> pairVector = vec.Vector<pair.Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair.Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

/*const unsigned int vertexCount = 2;

f<int> main() {
    /*int[vertexCount][vertexCount] graph = {
        { 0, 4, 0, 0, 0, 0, 0, 8, 0 },
        { 4, 0, 8, 0, 0, 0, 0, 11, 0 },
        { 0, 8, 0, 7, 0, 4, 0, 0, 2 },
        { 0, 0, 7, 0, 9, 14, 0, 0, 0 },
        { 0, 0, 0, 9, 0, 10, 0, 0, 0 },
        { 0, 0, 4, 14, 10, 0, 2, 0, 0 },
        { 0, 0, 0, 0, 0, 2, 0, 1, 6 },
        { 8, 11, 0, 0, 0, 0, 1, 0, 7 },
        { 0, 0, 2, 0, 0, 0, 6, 7, 0 }
    };

    printf("Test: %d\n", graph[1][7]);*/

    //int[vertexCount][5] graph = {{ 1, 2 }, { 3, 4 }, { 5, 6 }, { 7, 8 }, { 9, 10 }};
    /*unsafe {
        printf("Address: %p\n", &(*(&graph[2] + 0))[0]);
        printf("Value: %d\n", (*(&graph[2] + 0))[0]);
    }*/
    //printf("Result: %d\n", graph[2][1]);
    /*int[vertexCount][vertexCount] graph = {{ 1, 2 }, { 3, 4 }};
    int[vertexCount] graph1 = graph[0];
    printf("Test: %d\n", graph1[0]);
}*/

type T dyn;

f<int> main() {
    printf("Size: %d", sizeof(T));
}