import "std/text/analysis";

// Generic type definitions
type StrTy String|string;

// Prints the given string to the console
public inline p print<StrTy>(StrTy text) {
    printf("%s", text);
}

// Prints the given string to the console with a trailing line break
public inline p println<StrTy>(StrTy text) {
    printf("%s\n", text);
}

// Prints one or several line breaks to the console
public inline p lineBreak(unsigned int number = 1) {
    for int i = 0; i < number; i++ {
        printf("\n");
    }
}

public inline p beep() {
    printf("\a");
}

public p printColumn(string text, unsigned int width) {
    const unsigned long length = len(text);
    unsigned long i = 0l;

    while (i < length) {
        // Find the last word that fits within the width
        unsigned long j = i + width;
        while (j > i & j < length && !isWhitespace(text[j])) {
            j--;
        }
        // Print the word
        for (unsigned long k = i; k < j & k < length; k++) {
            printf("%c", text[k]);
        }
        // Move to the next line
        printf("\n");
        // Move to the next word
        i = j;
        while (i < length && isWhitespace(text[i])) {
            i++;
        }
    }
}

public p printColumn(const String& text, unsigned int width) {
    return this.printColumn(text.getRaw(), width);
}

public p printFixedWidth(string text, unsigned int width, bool ellipsis = false) {
    unsigned long length = len(text);
    const bool printEllipsis = ellipsis & length > width;

    for (unsigned long i = 0l; i < width; i++) {
        if (i < (printEllipsis ? cast<unsigned long>(width) - 3ul : length)) {
            printf("%c", text[i]);
        } else if (printEllipsis) {
            printf("...");
            break;
        } else {
            printf(" ");
        }
    }
}

public p printFixedWidth(const String& text, unsigned int width, bool ellipsis = false) {
    return this.printFixedWidth(text.getRaw(), width, ellipsis);
}
