type Test struct {
    double field1
    bool field2
}

f<byte> Test.getByte() {
    result = (byte) 12;
}

f<int> main() {
    dyn test = Test { 4.51, false };
    result = test.getInt();
}