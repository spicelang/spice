import "source1";

type Outer struct {
    int i
}

f<int> main() {
    TestStruct<Outer> _ts = TestStruct<Outer>();
}