/*import "std/data/vector" as vec;
import "std/data/pair" as pair;

f<int> main() {
    vec.Vector<pair.Pair<int, string>> pairVector = vec.Vector<pair.Pair<int, string>>();
    pairVector.pushBack(pair.Pair<int, string>(0, "Hello"));
    pairVector.pushBack(pair.Pair<int, string>(1, "World"));

    pair.Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!", p1.getSecond());
}*/

f<int> getAge() {
    dyn i;
    if (true) {
        result = 20;
        return;
    } else if (i = false) {
        result = 19;
    }
    return 15;
}

f<int> main() {
    int age = getAge();
    printf("The age is: %d", age);
}