f<int> main() {
    printf("Test");
}