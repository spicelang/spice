f<string> unusedFunction() {
    return "Test";
}

f<int> main() {}