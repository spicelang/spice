type Visitor struct {}

type SymbolTable struct {}

type Visitable interface {
    f<bool> accept(Visitor*);
}

type AstNode struct : Visitable {}

type AstEntryNode struct : Visitable {
    AstNode astNode
    SymbolTable* extFunctionScope
    bool takesArgs
}

f<int> main() {
    dyn entryNode = AstEntryNode{};
    printf("%d", entryNode.takesArgs);
}