#![core.compiler.alwaysKeepOnNameCollision = true]

// Link external functions
ext f<heap byte*> malloc(unsigned long);
ext f<heap byte*> realloc(heap byte*, unsigned long);
ext p free(heap byte*);
ext p memcpy(heap byte*, heap byte*, unsigned long);

// Generic type defs
type T dyn;

/**
  * Allocates a new block of memory of the given size.
  *
  * @param size The size of the block to allocate.
  * @return A pointer to the allocated block, or an error if the allocation failed.
  */
public f<Result<heap byte*>> sAlloc(unsigned long size) {
    heap byte* ptr = malloc(size);
    return ptr != nil<heap byte*> ? ok(ptr) : err<heap byte*>("Out of memory occurred!");
}

/**
  * Reallocates a block of memory to the given size.
  *
  * @param ptr The pointer to the block to reallocate.
  * @param size The new size of the block.
  * @return A pointer to the reallocated block, or an error if the reallocation failed.
  */
public f<Result<heap byte*>> sRealloc(heap byte* ptr, unsigned long size) {
    heap byte* newPtr = realloc(ptr, size);
    return newPtr != nil<heap byte*> ? ok(newPtr) : err<heap byte*>("Out of memory occurred!");
}

/**
  * Copies a block of memory to a new block of memory.
  *
  * @param oldPtr The pointer to the block to copy.
  * @param newPtr The pointer to the new block to copy to.
  * @param size The size of the block to copy.
  * @return A pointer to the copied block, or an error if the copy failed.
  */
public f<Result<heap byte*>> sCopy(heap byte* oldPtr, heap byte* newPtr, unsigned long size) {
    if oldPtr == nil<heap byte*> | newPtr == nil<heap byte*> {
        return err<heap byte*>("Cannot copy from or to nil pointer!");
    }
    memcpy(newPtr, oldPtr, size);
    return ok(newPtr);
}

/**
  * Frees a block of memory.
  * The pointer is zeroed out after freeing the memory to prevent accidental double frees.
  *
  * @param ptr The pointer to the block to free.
  */
public p sDealloc(heap byte*& ptr) {
    if ptr == nil<heap byte*> { return; }
    free(ptr);
    ptr = nil<heap byte*>; // Zero out to prevent accidental double frees
}

/**
 * Allocates memory for a new instance of the given type on the heap.
 * Note: This function panics if the allocation fails.
 *
 * @return A pointer to the heap-allocated instance
 */
public f<heap T*> sNew<T>() {
    unsafe {
        // Allocate memory for the instance
        Result<heap byte*> res = sAlloc(sizeof(type T));
        return (heap T*) res.unwrap();
    }
}

/**
 * Allocates memory for a new instance of the given type on the heap.
 * Note: This function panics if the allocation fails.
 *
 * @param val The value to put into the heap-allocated memory
 * @return A pointer to the heap-allocated instance
 */
public f<heap T*> sNew<T>(const T& val) {
    unsafe {
        // Allocate memory for the instance
        Result<heap byte*> res = sAlloc(sizeof(type T));
        result = (heap T*) res.unwrap();
        // Copy the value into the heap-allocated memory
        sCopy((heap byte*) &val, (heap byte*) result, sizeof(type T));
    }
}

/**
 * Allocates memory for a new instance of the given type on the heap.
 *
 * @param ptr The pointer to the heap-allocated memory
 * @param val The value to put into the heap-allocated memory
 * @return A pointer to the heap-allocated instance
 */
public f<T*> sPlacementNew<T>(heap byte* ptr, const T& val) {
    unsafe {
        // Copy the value into the heap-allocated memory
        sCopy((heap byte*) &val, ptr, sizeof(type T));
        return (T*) ptr;
    }
}

/**
 * Destroys the given heap-allocated instance and frees the memory.
 *
 * @param ptr The pointer to the heap-allocated instance
 */
public p sDelete<T>(heap T*& ptr) {
    unsafe {
        // Destruct the object
        ptr.dtor();
        // Deallocate the memory
        sDealloc((heap byte*&) ptr);
    }
}

/**
 * Creates a non-owned pointer to the given heap-allocated instance.
 *
 * @param ptr The pointer to the heap-allocated instance
 * @return A non-owned pointer to the heap-allocated instance
 */
public f<T*> sNonOwned<T>(heap T* ptr) {
    unsafe {
        return ptr;
    }
}
