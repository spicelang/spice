import "std/io/logging";
import "std/io/filepath";

f<int> main() {
    LogFile logFile = LogFile(FilePath("test.txt"), false);
    logFile.logDebug("This is a debug message");
    logFile.logInfo("This is a info message");
    logFile.logWarning("This is a warning message");
    logFile.logError("This is a error message");
}