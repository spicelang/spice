/*f<int> test(string input) {
    return 12;
}

p invoke(f<int>(string) fctPtr) {
    fctPtr("string");
}*/

f<int> test() {
    printf("Hi");
    return 12;
}

f<int> main() {
    int t = test();
    //f<int>(string) testFct = test;
    //invoke(testFct);
}