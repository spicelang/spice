f<int> main() {
    String strA = String("Hello ");
    String strB = String("World!");
    String strC = strA + strB;
    printf("%s\n", strA);
    printf("%s\n", strB);
    printf("%s\n", strC);
}