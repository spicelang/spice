// Prints the given string to the console
public p print(string text) {
    printf("%s", text);
}

// Prints the given string to the console with a trailing line break
public p println(string text) {
    printf("%s\n", text);
}

// Prints one or several line breaks to the console
public p lineBreak(unsigned int number = 1) {
    for int i = 0; i < number; i++ {
        printf("\n");
    }
}

public p beep() {
    printf("\a");
}