type TestStruct struct {
    int a
}

p TestStruct.unusedProcedure() {
    printf("Hello World: %d", this.a);
}

f<string> TestStruct.unusedFunction() {
    printf("%d", this.a);
    return "Hello World";
}

f<int> main() {
    TestStruct _ts;
}

/*type Parent struct {
    int i
}

type Child struct {
    compose Parent parent
    int j
    int k
}

f<int> main() {
    Child child;
    child.i = 3;
    child.j = 5;
}*/

/*import "std/os/env";
import "std/io/filepath";
import "bootstrap/ast/ast-nodes";
import "bootstrap/lexer/lexer";
import "bootstrap/parser/parser";

f<int> main() {
    String filePathString = getEnv("SPICE_STD_DIR") + "/../test/test-files/bootstrap-compiler/standalone-parser-test/test-file.spice";
    FilePath filePath = FilePath(filePathString);
    Lexer lexer = Lexer(filePath);
    Parser parser = Parser(lexer);
    ASTEntryNode* ast = parser.parse();
    assert ast != nil<ASTEntryNode*>;
    printf("All assertions passed!\n");
}*/