type T int|long;

type TestStruct<T> struct {
    unsigned T f1
    unsigned long length
}

f<int> main() {
    dyn a = TestStruct<long>{(unsigned long) 12345l, (unsigned long) 54321l};
}