//import "../../src-bootstrap/util/CodeLoc";
//import "../../src-bootstrap/ast/ASTNodes";

f<int> main() {
    //CodeLoc cl = CodeLoc(1l, 2l, "File path");
    //ASTNode node = ASTNode(nil<ASTNode*>, cl);
    dyn s4 = String("Hello World!");
    printf("%d", s4.rfind("o", 6l));
}