// Link external functions
ext f<byte*> malloc(long);
ext p free(byte*);

// Add generic type definitions
type T dyn;

/**
 * Node of a LinkedList
 */
public type Node<T> struct {
    T value
    Node<T>* next
}

/**
 * A linked list is a common, dynamically resizable data structure to store uniform data in order.
 * It is characterized by the pointer for each item, pointing to the next one.
 *
 * E.g. for a LinkedList<int>:
 * 1234 -> 4567 -> 7890 -> 4567 -> nil<int*>
 * tail                    head
 *
 * Time complexity:
 * Insert: O(1)
 * Delete: O(1)
 * Search: O(n)
 *
 * Beware that each add operation allocates memory and every remove operation frees memory.
 */
public type LinkedList<T> struct {
    Node<T>* tail
    Node<T>* head
}

public p LinkedList.ctor() {
    this.tail = nil<Node<T>*>;
    this.head = nil<Node<T>*>;
}

public p LinkedList.dtor() {
    Node<T>* curr = this.tail;
    while curr != nil<Node<T>*> {
        Node<T>* next = curr.next;
        free(curr);
        curr = next;
    }
}

public p LinkedList.insert(const T& value) {
    // Create new node
    Node<T>* newNode;
    unsafe {
        newNode = (Node<T>*) malloc(sizeof(type Node<T>) / 8l);
    }
    newNode.value = value;
    newNode.next = nil<Node<T>*>;

    // Insert at head
    this.head.next = newNode;
    this.head = newNode;
}

public p LinkedList.insertAt(unsigned long idx, const T& value) {
    // Create new node
    Node<T>* newNode;
    unsafe {
        newNode = (Node<T>*) malloc(sizeof(type Node<T>) / 8);
    }
    newNode.value = value;

    // Search for item right before insert position
    Node<T>* prev = this.tail;
    while curr != nil<Node<T>*> && idx > 1 {
        prev = prev.next;
        idx--;
    }

    // Link the next node to the new one
    newNode.next = prev.next;
    // Link the new node to the previous one
    prev.next = newNode;

    // Check if we have a new tail
    if idx == 0l {
        this.tail = newNode;
    }
    // Check if the previous node was the last node
    if this.head == prev {
        this.head = newNode;
    }
}

public p LinkedList.remove(const T& valueToRemove) {
    Node<T>* curr = this.tail;
    Node<T>* prev = nil<T*>;
    while curr != nil<Node<T>*> && curr.value != valueToRemove {
        prev = curr;
        curr = curr.next;
    }
    // Check if the item was found. If yes, delete its node
    if curr != nil<Node<T>*> {
        // Set the next node of the previous node
        prev.next = curr.next;
        // Free the removed node
        free(curr);
    }
}

public inline f<T&> LinkedList.getFirst() {
    return this.head.value;
}

public inline f<T&> LinkedList.getLast() {
    return this.tail.value;
}