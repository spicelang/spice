import "std/io/cli-subcommand";

// Generic types
type T bool|string|int|long|short;

public type CliParser struct {
    CliSubcommand rootSubcommand
}

public p CliParser.ctor(string appName, string appDescription = "") {
    this.rootSubcommand = CliSubcommand(nil<CliSubcommand*>, "v0.1.0", appName, appDescription);
}

public p CliParser.setVersion(string versionString) {
    this.rootSubcommand.setVersion(versionString);
}

public p CliParser.setFooter(string footer) {
    this.rootSubcommand.setFooter(footer);
}

public p CliParser.setRootCallback(p() callback) {
    this.rootSubcommand.setCallback(callback);
}

public p CliParser.allowUnknownOptions() {
    this.rootSubcommand.allowUnknownOptions();
}

public f<CliSubcommand&> CliParser.addSubcommand(string name, string description) {
    return this.rootSubcommand.addSubcommand(name, description);
}

public p CliParser.addOption<T>(string name, T& targetVariable, string description) {
    this.rootSubcommand.addOption(targetVariable, description);
}

public p CliParser.addFlag(string name, bool& targetVariable, string description) {
    this.rootSubcommand.addFlag(name, targetVariable, description);
}

public p CliParser.addFlag(string name, p(bool&) callback, string description) {
    this.rootSubcommand.addFlag(name, callback, description);
}

public f<int> CliParser.parse(unsigned int argc, string[] argv) {
    return this.rootSubcommand.parse(argc, argv);
}