f<int> main() {
    double doubleValue = 4.5;
    printf("Size: %d", sizeof(type doubleValue));
}