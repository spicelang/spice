f<int> main() {
    printf("Working ...");
    return 0;
    printf("Unreachable");
}