type Size alias long;

f<int> main() {
    printf("Do something different");
}