import "source1" as s1;
import "source2" as s2;

f<int> dummy() {
    return s1::dummy() + s2::dummy();
}

f<int> main() {
    int _res = dummy();
}