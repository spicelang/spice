import "std/io/file" as file;

f<int> main() {
    // Write to file
    file.writeFile("./test.txt", "Hello World\nThis is a test");
}