/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/net/socket" as socket;

f<int> main() {
    socket.Socket s = socket.openServerSocket(8080s, 2);
    printf("Error code: %d", s.errorCode);
    //s.close();
}*/


import "std/time/delay" as delay;

f<int> main() {
    int t1;
    int t2;
    int t3;

    t1 = thread {
        delay.delay(100);
        printf("Thread 1: %d, %d\n", tid(), t1);
        //join(t2);
        delay.delay(300);
        printf("Thread 1 finished\n");
    };

    t2 = thread {
        delay.delay(100);
        printf("Thread 2: %d, %d\n", tid(), t2);
        printf("tid(t1): %d\n", t1);
        printf("tid(t3): %d\n", t3);
        join(t1);
        printf("Thread 2 finished\n");
    };

    t3 = thread {
        delay.delay(100);
        printf("Thread 3: %d, %d\n", tid(), t3);
        delay.delay(200);
        printf("Thread 3 finished\n");
    };

    delay.delay(1000);
}