type StructToCopy struct {
    int a = 21
    bool b = false
}

f<int> main() {
    StructToCopy stc;
    printf("%d %d\n", stc.a, stc.b);
    StructToCopy stc2 = stc;
    printf("%d %d\n", stc2.a, stc2.b);
}