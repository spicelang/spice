import "std/os/dir" as dir;

f<int> main() {
    dir.createDir("./test.txt");
}