type Test struct {
    int i
    string s = "test"
}

f<int> main() {
    Test t;
    printf("Int: %d\n", t.i);
    printf("String: %s\n", t.s);
}

/*import "std/data/hash-table";

f<int> main() {
    HashTable<int, int> ht;
    ht.insert(1, 2);
    ht.insert(2, 3);
    ht.insert(3, 4);
    ht.insert(4, 5);
    ht.insert(5, 6);
}*/