import "source1";
import "source1";

f<int> main() {}