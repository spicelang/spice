// External declarations
ext f<long> strtol(string, char**, int);
ext f<int> atoi(string, char**, int);
ext f<double> strtod(string, char**);

// Converts a string to a double
public f<double> toDouble(string input) {
    return strtod(input, nil<char**>);
}

// Converts a string to an int
public f<int> toInt(string input, int base = 10) {
    return atoi(input, nil<char**>, base);
}

// Converts a string to a short
public f<short> toShort(string input, int base = 10) {
    return (short) atoi(input, nil<char**>, base);
}

// Converts a string to a long
public f<long> toLong(string input, int base = 10) {
    return strtol(input, nil<char**>, base);
}

// Converts a string to a byte
public f<byte> toByte(string input, int base = 10) {
    return (byte) atoi(input, nil<char**>, base);
}

// Converts a string to a char
public f<char> toChar(string input) {
    return input[0];
}

// Converts a string to a bool
public f<bool> toBool(string input) {
    return input == "true";
}