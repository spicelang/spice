// Link external functions
ext f<heap byte*> malloc(long);
ext p free(heap byte*);

// Add generic type definitions
type T dyn;

/**
 * Node of a BinaryTree
 */
public type Node<T> struct {
    heap Node<T>* childLeft
    heap Node<T>* childRight
    T value
}

/**
 * A binary tree is a data structure to fasten up search speeds. Binary trees (when balanced) can be searched in O(log n).
 * Insert operations, on the other hand, are rather slow, because the tree might get re-balanced.
 *
 * Time complexity:
 * Insert: O(n * m); n = inserted elements, m = moved elements
 * Delete: O(n * m); n = deleted elements, m = moved elements
 * Search: O(log n)
 */
public type BinaryTree<T> struct {
    heap Node<T>* rootNode
    bool isBalanced
}

public p BinaryTree.ctor() {
    this.rootNode = nil<heap Node<T>*>;
    this.isBalanced = false;
}

public p BinaryTree.dtor() {
    if this.rootNode != nil<heap Node<T>*> {
        this.rootNode.dtor();
        free((heap byte*) this.rootNode);
    }
}

public p Node.dtor() {
    if this.childLeft != nil<heap Node<T>*> {
        this.childLeft.dtor();
        free((heap byte*) this.childLeft);
    }
    if this.childRight != nil<heap Node<T>*> {
        this.childRight.dtor();
        free((heap byte*) this.childRight);
    }
}

public p BinaryTree.insert<T>(T newValue, heap Node<T>* baseNode = nil<heap Node<T>*>) {
    // Search position where to insert
    // ToDo
}