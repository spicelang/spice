f<double> testFunction(double param1) {
    result = 4.1;
}

f<int> main() {
    testFunction();
}