import "std/type/any";

public type AbstractAstVisitor interface {
    f<Any> visitEntry(EntryNode*);
    f<Any> visitMainFctDef(EntryNode*);
    f<Any> visitFctDef(EntryNode*);
    f<Any> visitProcDef(EntryNode*);
}