// Constants
const unsigned int INITIAL_ALLOC_COUNT = 5;
const unsigned int RESIZE_FACTOR = 2;

// Link external functions
ext<char*> malloc(int);
ext free(char*);
ext<char*> memcpy(char*, char*, int);

// Add generic type definition
type T dyn;

/**
 * A vector in Spice is a commonly used data structure, which can be used to represent a list of items
 */
public type Vector<T> struct {
    T* contents             // Pointer to the first data element
    unsigned long capacity  // Allocated number of items
    unsigned long size      // Current number of items
    unsigned int itemSize   // Size of a single item
}

public p Vector.constructor() {
    // Allocate space for the initial number of elements
    this.itemSize = sizeof(*this.contents);
    this.contents = malloc(this.itemSize * INITIAL_ALLOC_COUNT);
    this.capacity = INITIAL_ALLOC_COUNT;
}

public p Vector.destructor() {
    // Free all the memory
    free(this.contents);
}

/**
 * Add an item at the end of the vector
 */
public p Vector.pushBack<T>(T item) {
    // Check if we need to re-allocate memory
    if this.isFull() {
        this.capacity *= RESIZE_FACTOR;
        this.contents = malloc(this.itemSize * this.capacity);
    }

    // Insert the element at the back
    this.contents[this.size++] = item;
}

/**
 * Removes all items from the vector
 */
public p Vector.clear() {
    this.size = 0;
}

/**
 * Retrieve the current size of the queue
 *
 * @return Current size of the queue
 */
public f<long> Vector.size() {
    return this.size;
}

/**
 * Checks if the queue contains any items at the moment
 *
 * @return Empty or not empty
 */
public f<bool> Vector.isEmpty() {
    return this.size == 0l;
}

/**
 * Checks if the queue exhausts its capacity and needs to resize at the next call of push
 *
 * @return Full or not full
 */
public f<bool> Vector.isFull() {
    return this.size == this.capacity;
}

/**
 * Frees allocated memory that is not used by the queue
 */
public p Vector.pack() {
    // Return if no packing is required
    if this.isFull() { return; }
    // Pack the array
    this.resize(this.size);
}

/**
 * Re-allocates heap space for the queue contents
 */
p Vector.resize(unsigned long itemCount) {
    // Allocate the new memory
    T* newMemory = malloc(this.itemSize * itemCount);
    // Copy contents over
    memcpy(newMemory, this.contents, this.itemSize * this.capacity);
    // Free the old memory
    free(this.contents);
    // Set new memory to contents array
    this.contents = newMemory;
    this.capacity = itemCount;
}