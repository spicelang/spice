type TestStruct struct {
    int value
    len int
}

f<int> main() {
    printf("Test");
}