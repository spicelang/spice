import "test3" as s3;

public f<int> dummy() {
    return 1;
}