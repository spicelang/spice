type A dyn;

p printFormat<A>(A element) {
    printf("Sizeof output: %d\n", sizeof(element));
}