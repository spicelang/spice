// Contains the operating system name in lower case
public const string OS_NAME = "linux";

// Contains the native path separator
public const char PATH_SEPARATOR = '/';

// Returns if the current OS is Linux
public f<bool> isLinux() {
    return true;
}

// Returns if the current OS is Windows
public f<bool> isWindows() {
    return false;
}