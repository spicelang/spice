// Std imports
import "std/text/print";
import "std/data/pair";
import "std/data/unordered-map";
import "std/data/vector";
import "std/io/filepath";

// Own imports
import "bootstrap/driver";
//import "bootstrap/global/global-resource-manager";
import "bootstrap/ast/ast-nodes";
import "bootstrap/bindings/llvm/llvm";
import "bootstrap/util/compiler-warning";
import "bootstrap/symboltablebuilder/symbol-table-entry";
import "bootstrap/symboltablebuilder/scope";

type CompileStageType enum {
    NONE,
    LEXER,
    PARSER,
    CST_VISUALIZER,
    AST_BUILDER,
    AST_VISUALIZER,
    IMPORT_COLLECTOR,
    SYMBOL_TABLE_BUILDER,
    TYPE_CHECKER_PRE,
    TYPE_CHECKER_POST,
    IR_GENERATOR,
    IR_OPTIMIZER,
    OBJECT_EMITTER,
    FINISHED
}

type CompileStageIOType enum {
    IO_CODE,
    IO_TOKENS,
    IO_CST,
    IO_AST,
    IO_IR,
    IO_OBJECT_FILE
}

type TimerOutput struct {
  unsigned long lexer = 0l
  unsigned long parser = 0l
  unsigned long cstVisualizer = 0l
  unsigned long astBuilder = 0l
  unsigned long astVisualizer = 0l
  unsigned long importCollector = 0l
  unsigned long symbolTableBuilder = 0l
  unsigned long typeCheckerPre = 0l
  unsigned long typeCheckerPost = 0l
  unsigned long irGenerator = 0l
  unsigned long irOptimizer = 0l
  unsigned long objectEmitter = 0l
}

/**
 * Collects the output of the compiler for debugging
 */
type CompilerOutput struct {
    String cstString
    String astString
    String symbolTableString
    String irString
    String irOptString
    String asmString
    String typesString
    Vector<CompilerWarning> warnings
    TimerOutput times
}

type NameRegistryEntry struct {
    String name
    unsigned long typeId // Set for structs, interfaces and enums
    SymbolTableEntry* targetEntry
    Scope* targetScope
    SymbolTableEntry* importEntry = nil<SymbolTableEntry*>
}

/**
 * Represents a single source file
 */
public type SourceFile struct {
    // Public fields
    public String name
    public String fileName
    public FilePath filePath
    public String fileDir
    public bool isStdFile = false
    public bool isMainFile = true
    public bool alwaysKeepSymbolsOnNameCollision = false
    public bool ignoreWarnings = false
    public CompileStageType previousStage = CompileStageType::NONE
    public CompilerOutput compilerOutput
    public SourceFile* parent
    public String cacheKey
    public bool restoredFromCache = false
    public EntryNode* ast = nil<EntryNode*>
    public heap Scope* globalScope
    public llvm::LLVMContext context
    public llvm::IRBuilder builder
    public heap llvm::TargetMachine* targetMachine
    public heap llvm::Module* llvmModule
    public UnorderedMap<String, SourceFile*> dependencies
    public Vector<const SourceFile*> dependants
    public Map<String, NameRegistryEntry> exportedNameRegistry
    public Vector<const Function*> testFunctions
    // Private fields
    GlobalResourceManager& resourceManager
    CliOptions& cliOptions
    UnorderedMap<const Type*, llvm::Type*> llvmTypeMapping
    unsigned short importedRuntimeModules = 0s
    unsigned short totalTypeCheckerRuns = 0s
}

public p SourceFile.ctor(GlobalResourceManager &resourceManager, SourceFile* parent, const String& name, const String& filePath, bool isStdFile) {
    // Copy data
    this.resourceManager = resourceManager;
    this.parent = parent;
    this.name = name;
    this.filePath = filePath;
    this.isStdFile = isStdFile;

    // Deduce fileName and fileDir
    /*this.fileName = ;
    this.fileDir = ;*/
}

public p SourceFile.runLexer() {
    // Lex this source file
}

public p SourceFile.runParser() {
    // Parse this source file
}

public p SourceFile.runCSTVisualizer(string* output) {
    // Only execute if enabled
    if !cliOptions.dumpCST && !cliOptions.testMode { return; }

    // ToDo: Extend
}

public p SourceFile.runASTBuilder() {
    // Transform the imported source files
    // ToDo: Extend
}

public p SourceFile.runASTVisualizer(string* output) {
    // Only execute if enabled
    if !cliOptions.dumpAST && !cliOptions.testMode { return; }

    // ToDo: Extend
}

public p SourceFile.runImportCollector() {

}

public p SourceFile.runSymbolTableBuilder() {

}

public p SourceFile.runTypeChecker() {

}

p SourceFile.runTypeCheckerPre() {

}

p SourceFile.runTypeCheckerPost() {

}

public p SourceFile.runIRGenerator() {

}

public p SourceFile.runDefaultIROptimizer() {

}

public p SourceFile.runObjectEmitter() {

}

public p SourceFile.concludeCompilation() {

}

public p SourceFile.runFrontEnd() {

}

public p SourceFile.runMiddleEnd() {

}

public p SourceFile.runBackEnd() {

}

f<bool> SourceFile.isAlreadyImported(const String& filePathSearch) {
    // Check if the current source file corresponds to the path to search
    if this.filePath == filePathSearch { return true; }
    // Check parent recursively
    return this.parent != nil<SourceFile*> && this.parent.isAlreadyImported(filePathSearch);
}