import "std/data/stack" as s;

f<int> main() {
    dyn doubleVec = s.Stack<double>(3, 6.4);
    printf("Test: %f\n", doubleVec.pop());
    printf("Test: %f\n", doubleVec.pop());
    printf("Test: %f\n", doubleVec.pop());
    printf("Test: %f\n", doubleVec.pop());
    doubleVec.dtor();
}