#![core.compiler.alwaysKeepOnNameCollision = true]

/**
 * This is the generalized error type in Spice and part of the error handling mechanism.
 */
public type Error struct {
    public int code
    public string message
}

public p Error.ctor() {
    this.code = 0;
    this.message = "Runtime error";
}

public p Error.ctor(int errorCode, string message) {
    this.code = errorCode;
    this.message = message;
}

public p Error.ctor(string message) {
    this.code = 1;
    this.message = message;
}

/**
 * Prints the error message to the console.
 */
public p Error.print() {
    printf("%s\n", this.message);
}

/**
 * Panic with this error
 */
public p Error.toPanic() {
    panic(*this);
}