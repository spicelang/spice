// Std imports
import "std/data/unordered-map";
import "std/data/vector";

// Own imports
import "bootstrap/ast/ast-nodes";
import "bootstrap/reader/code-loc";
import "bootstrap/symboltablebuilder/qual-type";
import "bootstrap/symboltablebuilder/scope-intf";
import "bootstrap/symboltablebuilder/symbol-table-entry";
import "bootstrap/symboltablebuilder/type-qualifiers";
import "bootstrap/symboltablebuilder/capture";
import "bootstrap/model/generic-type";
import "bootstrap/model/function";
import "bootstrap/model/struct";
import "bootstrap/model/interface";
import "bootstrap/util/compiler-warning";

// Type aliases
public type CaptureMap alias UnorderedMap</*name=*/string, /*capture*/Capture>;
public type SymbolMap alias UnorderedMap</*name=*/string, /*entry*/SymbolTableEntry>;

/**
 * Class for storing information about symbols of the program.
 * Symbol tables are arranged in a tree structure, so that you can navigate with the .parent property and getChild() method up
 * and down the tree.
 */
public type SymbolTable struct {
    SymbolTable* parent
    IScope* scope
    SymbolMap symbols
    CaptureMap captures
    bool capturingRequired = false
}

public p SymbolTable.ctor(SymbolTable* parent, IScope* scope) {
    this.parent = parent;
    this.scope = scope;
}

/**
 * Insert a new symbol into the current symbol table. If it is a parameter, append its name to the paramNames vector
 *
 * @param name Name of the symbol
 * @param declNode AST node where the symbol is declared
 * @return Inserted entry
 */
public p SymbolTable.insert(const String& name, const ASTNode* declNode) {
    const bool isGlobal = this.parent == nil<SymbolTable*>;
    const unsigned int orderIndex = this.symbols.getSize();
    // Insert into symbols map. The type is 'dyn', because concrete types are determined by the type checker later on
    // ToDo: Implement
}

/**
 * Insert a new anonymous symbol into the current symbol table.
 * The anonymous symbol will be identified via the definition code location
 *
 * @param qualType Type of the symbol
 * @param declNode AST node where the anonymous symbol is declared
 * @return Inserted entry
 */
public p SymbolTable.insertAnonymous(const QualType& qualType, ASTNode* declNode, unsigned long numericSuffix = 0l) {
    // ToDo: Implement
}

/**
 * Copy a symbol by its name
 *
 * @param originalName Original symbol name
 * @param newName New symbol name
 * @return Copied entry
 */
public f<SymbolTableEntry*> SymbolTable.copySymbol(const String& originalName, const String& newName) {
    SymbolTableEntry* entryToCopy = lookupStrict(originalName);
    assert entryToCopy != nil<SymbolTableEntry*>;
    // ToDo
    return nil<SymbolTableEntry*>;
}

/**
 * Check if a symbol exists in the current or any parent scope and return it if possible
 *
 * @param name Name of the desired symbol
 * @return Desired symbol / nullptr if the symbol was not found
 */
public f<SymbolTableEntry*> SymbolTable.lookup(const String& name) {
    // Check if the symbol exists in the current scope. If yes, take it
    SymbolTableEntry* entry = this.lookupStrict(name);
    if entry == nil<SymbolTableEntry*> { // Symbol was not found in the current scope
        // We reached the root scope, the symbol does not exist at all
        if parent == nil<SymbolTable*> {
            return nil<SymbolTableEntry*>;
        }
        // If there is a parent scope, continue the search there
        entry = this.parent.lookup(name);
        // Symbol was also not found in all the parent scopes, return nullptr
        if entry == nil<SymbolTable*> {
            return nil<SymbolTableEntry*>;
        }

        // Check if this scope requires capturing and capture the variable if appropriate
        const QualType entryType = entry.getQualType();
        if this.capturingRequired && !this.captures.contains(name) && !entryType.isOneOf([TY_IMPORT, TYPE_FUNCTION, TY_PROCEDURE]) {
            // We need to make the symbol volatile if we are in an async scope and try to access a symbol that is not in an async scope
            entry.isVolatile = this.scope.isInAsyncScope() && !entry.scope.isInAsyncScope();
            // Add the capture to the current scope
            this.captures.insert(name, Capture(entry));
        }
    }
    return entry;
}

/**
 * Check if a symbol exists in the current scope and return it if possible
 *
 * @param name Name of the desired symbol
 * @return Desired symbol / nullptr if the symbol was not found
 */
public f<SymbolTableEntry*> SymbolTable.lookupStrict(const string name) {
    if name.isEmpty() {
        return nil<SymbolTableEntry*>;
    }
    // Check if a symbol with this name exists in this scope
    if this.symbols.contains(name) {
        return &this.symbols.get(name);
    }
    // Check if a capture with this name exists in this scope
    if this.captures.contains(name) {
        return &this.captures.get(name).capturedSymbol;
    }
    // Otherwise, return a nullptr
    return nil<SymbolTableEntry*>;
}

/**
 * Check if a symbol exists in one of the composed field scopes of the current scope and return it if possible.
 * This only works if the current scope is a struct scope.
 *
 * @param name Name of the desired symbol
 * @param indexPath How to index the found symbol using order indices (e.g. for GEP)
 * @return Desired symbol / nullptr if the symbol was not found
 */
public f<SymbolTableEntry*> SymbolTable.lookupInComposedFields(const String& name, Vector<unsigned long> indexPath) {
    assert this.scopeType == ScopeType::STRUCT;
    // ToDo

    // Symbol was not found in current scope, return nullptr
    return nil<SymbolTableEntry*>;
}

/**
 * Check if an order index exists in the current or any parent scope and returns it if possible.
 * Warning: Unlike the `lookup` method, this one doesn't consider the parent scopes
 *
 * @param orderIndex Order index of the desired symbol
 * @return Desired symbol / nullptr if the symbol was not found
 */
public f<SymbolTableEntry*> SymbolTable.lookupStrictByIndex(const unsigned int orderIndex) {
    // ToDo
    return nil<SymbolTableEntry*>;
}

/**
 * Check if an anonymous symbol exists in the current scope and return it if possible
 *
 * @param codeLoc Definition code loc
 * @param numericSuffix Numeric suffix of the anonymous symbol
 * @return Anonymous symbol
 */
public f<SymbolTableEntry*> SymbolTable.lookupAnonymous(const CodeLoc& codeLoc) {
    const String name = String("anon.") + codeLoc.toString();
    if numericSuffix > 0 {
        name += '.';
        name += toString(numericSuffix);
    }
    return this.lookup(name);
}

/**
 * Check if a capture exists in the current or any parent scope scope and return it if possible
 *
 * @param name Name of the desired captured symbol
 * @return Capture / nullptr if the capture was not found
 */
public f<Capture> SymbolTable.lookupCapture(const String& name) {
    // Check if the capture exists in the current scope. If yes, take it
    Capture* capture = this.lookupCaptureStrict(name);
    if capture != nil<Capture*> {
        return capture;
    }

    // We reached the root scope, the symbol does not exist at all
    if this.parent == nil<SymbolTable*> {
        return nullptr;
    }

    return this.parent.lookupCapture(name);
}

/**
 * Check if a capture exists in the current scope and return it if possible
 *
 * @param name Name of the desired captured symbol
 * @return Capture / nullptr if the capture was not found
 */
public f<Capture> SymbolTable.lookupCaptureStrict(const string captureName) {
    // If available in the current scope, return it
    if this.captures.contains(captureName) {
        return &this.captures.get(captureName);
    }
    // Otherwise, return nullptr
    return nil<Capture*>;
}

/**
 * Set capturing for this scope to required.
 */
public p SymbolTable.setCapturingRequired() {
    this.capturingRequired = true;
}

/**
 * Deletes an existing anonymous symbol
 *
 * @param name Anonymous symbol name
 */
public p SymbolTable.deleteAnonymous(const String& name) {
    // ToDo
}

/**
 * Stringify a symbol table to a human-readable form. This is used to realize dumps of symbol tables
 *
 * Example:
 * {
 *   "name": "<SymbolTableName>"
 *   "symbols": [
 *     ... (SymbolTableEntry)
 *   ],
 *   "children": [
 *     ... (SymbolTable)
 *   ]
 * }
 *
 * @return Symbol table if form of a string
 */
public f<String> SymbolTable.toJSON() {
    // ToDo
    return String();
}
