import "std/data/unordered-map";

f<int> main() {
    UnorderedMap<int, string> map = UnorderedMap<int, string>(3l);
    assert map.getSize() == 0;
    assert map.isEmpty();
    map.upsert(1, "one");
    map.upsert(2, "two");
    map.upsert(3, "three");
    map.upsert(4, "four");
    assert map.getSize() == 4;
    assert !map.isEmpty();
    assert map.contains(1);
    assert map.contains(2);
    assert map.contains(3);
    assert map.contains(4);
    assert !map.contains(5);
    assert map.get(1) == "one";
    assert map.get(2) == "two";
    assert map.get(3) == "three";
    assert map.get(4) == "four";
    const Result<string> item5 = map.getSafe(5);
    assert item5.isErr();
    map.remove(2);
    assert !map.contains(2);
    assert map.getSize() == 3;
    map.clear();
    assert map.getSize() == 0;
    assert map.isEmpty();
    map.upsert(1, "one");
    map.upsert(1, "one new");
    assert map.getSize() == 1;
    assert map.get(1) == "one new";
    map.remove(1);
    assert map.isEmpty();

    printf("All assertions passed!\n");
}