//import "std/iterator/number-iterator";
import "std/runtime/iterator_rt";

f<int> main() {
    Vector<int> vi = Vector<int>();
    vi.pushBack(123);
    vi.pushBack(4321);
    dyn it = iterate(vi);
    printf("Get: %d\n", it.get());
    /*foreach int i : it {
        printf("Item: %d\n", i);
    }*/
}