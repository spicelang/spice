import "std/os/thread";

f<int> fib(int n) {
    if n <= 2 { return 1; }
    return fib(n - 1) + fib(n - 2);
}

f<int> main() {
    int threadCount = 8;
    Thread[8] threads = [];
    for unsigned int i = 0; i < threadCount; i++ {
        threads[i] = Thread(p() {
            int res = fib(30);
            printf("Thread returned with result: %d\n", res);
        });
        Thread& thread = threads[i];
        thread.run();
    }
    printf("Started all threads. Waiting for results ...\n");
    for unsigned int i = 0; i < threadCount; i++ {
        Thread& thread = threads[i];
        thread.join();
    }
    printf("Program finished");
}

/*import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

type ASTNode struct {
    int value
}

public p ASTNode.dtor() {
    printf("Dtor called!");
}

f<int> main() {
    DefaultMemoryManager defaultMemoryManager;
    IMemoryManager* memoryManager = &defaultMemoryManager;
    BlockAllocator<ASTNode> allocator = BlockAllocator<ASTNode>(memoryManager, 10l);
}*/