public const int SIZE = 64;
public const double MIN_VALUE = 0; // ToDo: Fix
public const double MAX_VALUE = 0; // ToDo: Fix

// Converts a double to an int
public f<int> toInt(double input) {
    // ToDo: Implement
    return 0;
}

// Converts a double to a short
public f<short> toInt(double input) {
    // ToDo: Implement
    return (short) 0;
}

// Converts a double to a long
public f<long> toInt(double input) {
    // ToDo: Implement
    return (long) 0;
}

// Converts a double to a byte
public f<byte> toByte(double input) {
    // ToDo: Implement
    result = (byte) 0;
}

// Converts a double to a string
public f<string> toString(double input) {
    // ToDo: Implement
    return "";
}

// Converts a double to a boolean
public f<bool> toBool(double input) {
    return input >= 0.5;
}