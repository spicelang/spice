import "std/os/env";

public f<string> getTempDir() {
    Result<string> dir = getEnv("TMPDIR");
    return dir.isOk() ? dir.unwrap() : "/tmp";
}
