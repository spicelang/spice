import "std/type/double" as doubleTy;

f<int> main() {
    // toInt()
    //int asInt = doubleTy.toInt(123.54);
    //assert asInt == 123;

    // toShort()
    //short asShort = doubleTy.toShort(12.345);
    //assert asShort == 12;

    // toLong()
    //long asLong = doubleTy.toLong(534569.2345);
    //assert asLong == 534569l;

    // toByte()
    //long asByte = doubleTy.toLong(53.89);
    //assert asByte == (byte) 53;

    // toString()
    //string asString = doubleTy.toString(9.0);
    //assert asString == "9.0";

    // toBool()
    bool asBool1 = doubleTy.toBool(1.0);
    assert asBool1 == true;
    bool asBool2 = doubleTy.toBool(0.0);
    assert asBool2 == false;

    printf("All assertions succeeded");
}