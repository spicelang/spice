f<int> main() {
    fallthrough;
}