import "std/type/type-conversion";

f<int> main() {
    // toDouble()
    double asDouble = toDouble("5.67");
    assert asDouble == 5.67;

    // toInt()
    int asInt = toInt("-6546");
    assert asInt == -6546;

    // toLong()
    long asLong = toLong("56");
    assert asLong == 56l;

    // toShort()
    short asShort = toShort("-12");
    assert asShort == -12s;

    // toByte()
    byte asByte = toByte("12");
    assert asByte == cast<byte>(12);

    // toChar()
    char asChar = toChar("i");
    assert asChar == 'i';

    // toBool()
    bool asBool1 = toBool("true");
    assert asBool1 == true;
    bool asBool2 = toBool("false");
    assert asBool2 == false;

    printf("All assertions succeeded");
}