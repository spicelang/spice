import "std/os/thread";
import "std/data/vector";
import "std/data/queue";
import "std/os/atomic";
import "std/os/cpu";
import "std/os/system";
import "std/runtime/iterator_rt";

/**
 * A thread pool that can be used to run multiple jobs in parallel.
 * Thread pools in Spice work with a fixed number of worker threads, that are created when the pool is started. After that, an
 * arbitrary number of jobs can be queued to be run by the pool. The pool will then run as many jobs as possible in parallel.
 */
public type ThreadPool struct {
    Vector<Thread> workerThreads
    Queue<p()> queuedJobs
    Atomic<unsigned short> runningJobs
    unsigned short workerThreadCount
    bool stopRequested = false
    bool stopOnEmptyQueueRequested = false
    bool pauseRequested = false
}

/**
 * Create a new thread pool.
 *
 * @param maxConcurrentJobs The maximum number of jobs that can be run at the same time. If 0, the number of CPU cores is used.
 */
public p ThreadPool.ctor(unsigned short workerThreadCount = 0s) {
    this.workerThreads = Vector<Thread>();
    this.queuedJobs = Queue<p()>();
    this.runningJobs = Atomic<unsigned short>(0s);
    this.workerThreadCount = workerThreadCount > 0s ? workerThreadCount : (unsigned short) getCPUCoreCount();
}

/**
 * Start the thread pool.
 */
public p ThreadPool.start() {
    p() workerRoutine = p() [[async]] {
        do {
            // Check if there are jobs to run
            const bool hasQueuedJobs = !this.queuedJobs.isEmpty();
            // If we are supposed to stop when the queue is empty and there are no more jobs, abort
            if this.stopOnEmptyQueueRequested & !hasQueuedJobs {
                break;
            }
            // If we are not supposed to stop and there are jobs, run them
            if !this.pauseRequested & hasQueuedJobs {
                p() task = this.queuedJobs.pop();
                this.runningJobs.store(this.runningJobs.load() + 1s);
                task();
                this.runningJobs.store(this.runningJobs.load() - 1s);
            }
            // Yield to other threads
            yield();
        } while (!this.stopRequested);
    };

    // Create worker threads
    for unsigned short i = 0s; i < this.workerThreadCount; i++ {
        this.workerThreads.pushBack(Thread(workerRoutine));
        Thread& workerThread = this.workerThreads.back();
        workerThread.run();
    }
    sizeof(0);
}

/**
 * Finish the running jobs and stop the thread pool.
 */
public p ThreadPool.stop() {
    // Stop worker threads
    this.stopRequested = true;
    // Wait for all worker threads to terminate
    this.joinWorkerThreads();
    // Reset the stop flag
    this.stopRequested = false;
}

/**
 * Wait for all queued jobs to finish and stop the thread pool.
 */
public p ThreadPool.join() {
    // Stop worker threads
    this.stopOnEmptyQueueRequested = true;
    // Wait for all worker threads to terminate
    this.joinWorkerThreads();
    // Reset the stop flag
    this.stopOnEmptyQueueRequested = false;
}

/**
 * Enqueue a job to be run by the thread pool.
 *
 * @param job The job routine to enqueue.
 */
public p ThreadPool.enqueue(const p()& job) {
    this.queuedJobs.push(job);
}

/**
 * Pause the thread pool. The worker threads will finish their current job and then wait for the pool to be resumed.
 */
public p ThreadPool.pause() {
    this.pauseRequested = true;
}

/**
 * Resume the thread pool.
 */
public p ThreadPool.resume() {
    this.pauseRequested = false;
}

/**
 * Check if the thread pool is paused.
 */
public f<bool> ThreadPool.isPaused() {
    return this.pauseRequested;
}

/**
 * Retrieve the number of jobs that are currently running.
 */
public f<unsigned short> ThreadPool.getRunningJobCount() {
    return this.runningJobs.load();
}

/**
 * Retrieve the number of jobs that are currently queued.
 */
public f<unsigned short> ThreadPool.getQueuedJobCount() {
    return (unsigned short) this.queuedJobs.getSize();
}

/**
 * Retrieve the number of worker threads.
 */
public f<unsigned short> ThreadPool.getWorkerThreadCount() {
    return this.workerThreadCount;
}

/**
 * Wait for all worker threads to terminate.
 */
p ThreadPool.joinWorkerThreads() {
    foreach const Thread& workerThread : this.workerThreads.getIterator() {
        workerThread.join();
    }
}