// Std imports
import "std/data/vector";
import "std/data/pair";

// Own imports
import "bootstrap/source-file-intf";
import "bootstrap/ast/ast-node-intf";
import "bootstrap/symboltablebuilder/super-type";
import "bootstrap/symboltablebuilder/type-intf";
import "bootstrap/symboltablebuilder/type-qualifiers";
import "bootstrap/symboltablebuilder/scope-intf";
import "bootstrap/model/function-intf";
import "bootstrap/model/struct-intf";
import "bootstrap/model/interface-intf";
import "bootstrap/model/generic-type-intf";

// Constants
public const string STROBJ_NAME = "String";
public const string RESULTOBJ_NAME = "Result";
public const string ERROBJ_NAME = "Error";
public const string TIOBJ_NAME = "TypeInfo";
public const string IITERATOR_NAME = "IIterator";
public const string ARRAY_ITERATOR_NAME = "ArrayIterator";
public const unsigned long TYPE_ID_ITERATOR_INTERFACE = 255ul;
public const unsigned long TYPE_ID_ITERABLE_INTERFACE = 256ul;

public type QualType struct {
    const IType* rawType = nil<const IType*>
    TypeQualifiers qualifiers
}

public type QualTypeList alias Vector<QualType>;
public type Arg alias Pair</*type=*/QualType, /*isTemporary=*/bool>;
public type ArgList alias Vector</*arg=*/Arg>;

public p QualType.ctor(SuperType superType) {

}

public p QualType.ctor(SuperType superType, const String& subType) {

}

public p QualType.ctor(const IType* rawType, TypeQualifiers qualifiers) {
    this.rawType = rawType;
    this.qualifiers = qualifiers;
}

/**
 * Get the super type of the underlying type
 *
 * @return Super type
 */
public f<SuperType> QualType.getSuperType() {
    return this.rawType.getSuperType();
}

/**
 * Get the subtype of the underlying type
 *
 * @return Subtype
 */
public f<const String&> QualType.getSubType() {
    return this.rawType.getSubType();
}

/**
 * Get the array size of the underlying type
 *
 * @return Array size
 */
public f<unsigned int> QualType.getArraySize() {
    return this.rawType.getArraySize();
}

/**
 * Get the body scope of the underlying type
 *
 * @return Body scope
 */
public f<IScope*> QualType.getBodyScope() {
    return this.rawType.getBodyScope();
}

/**
 * Get the function parameter types of the underlying type
 *
 * @return Function parameter types
 */
public f<QualType&> QualType.getFunctionReturnType() {
    return this.rawType.getFunctionReturnType();
}

/**
 * Get the function parameter types of the underlying type
 *
 * @return Function parameter types
 */
public f<QualTypeList> QualType.getFunctionParamTypes() {
    return this.rawType.getFunctionParamTypes();
}

/**
 * Get the function parameter and return types of the underlying type
 *
 * @return Function parameter and return types
 */
public f<QualTypeList&> QualType.getFunctionParamAndReturnTypes() {
    return this.rawType.getFunctionParamAndReturnTypes();
}

/**
 * Check if the underlying type has lambda captures
 *
 * @return Has lambda captures or not
 */
public f<bool> QualType.hasLambdaCaptures() {
    return this.rawType.hasLambdaCaptures();
}

/**
 * Get the template types of the underlying type
 *
 * @return Template types
 */
public f<QualTypeList&> QualType.getTemplateTypes() {
    return this.rawType.getTemplateTypes();
}

/**
 * Get the struct instance for a struct type
 *
 * @param node Accessing AST node
 * @return Struct instance
 */
public f<IStruct*> QualType.getStruct(const IASTNode* node) {
    assert this.is(SuperType::TY_STRUCT);
    IScope* structScope = this.getBodyScope();
    const String& structName = this.getSubType();
    const QualTypeList& templateTypes = this.getTemplateTypes();
    return matchStruct(structScope.getParent(), structName, templateTypes, node);
}

/**
 * Get the interface instance for an interface type
 *
 * @param node Accessing AST node
 * @return Interface instance
 */
public f<IInterface*> QualType.getInterface(const IASTNode* node) {
    assert this.is(SuperType::TY_INTERFACE);
    IScope* interfaceScope = this.getBodyScope();
    const String& interfaceName = this.getSubType();
    const QualTypeList& templateTypes = this.getTemplateTypes();
    return matchInterface(interfaceScope.getParent(), interfaceName, templateTypes, node);
}

/**
 * Check if the underlying type is of a certain super type
 *
 * @param superType Super type
 * @return Is of super type or not
 */
public f<bool> QualType.is(SuperType superType) {
    return this.rawType.is(superType);
}

/**
 * Check if the underlying type is one of a list of super types
 *
 * @param superTypes List of super types
 * @return Is one of the super types or not
 */
public f<bool> QualType.isOneOf(SuperType[] superTypes, unsigned long superTypesSize) {
    return this.rawType.isOneOf(superTypes, superTypesSize);
}

/**
 * Check if the base type of the underlying type is a certain super type
 *
 * @param superType Super type
 * @return Is base type or not
 */
public f<bool> QualType.isBase(SuperType superType) {
    return this.rawType.isBase(superType);
}

/**
 * Check if the underlying type is a primitive type
 * Note: enum types are mapped to int, so they are also count as primitive types.
 *
 * @return Primitive or not
 */
public f<bool> QualType.isPrimitive() {
    return this.rawType.isPrimitive();
}

/**
 * Check if the underlying type is an extended primitive type
 * The definition of extended primitive types contains all primitive types plus the following:
 * - structs
 * - interfaces
 * - functions/procedures
 *
 * @return Extended primitive or not
 */
public f<bool> QualType.isExtendedPrimitive() {
    return this.rawType.isExtendedPrimitive();
}

/**
 * Check if the underlying type is a pointer
 *
 * @return Pointer or not
 */
public f<bool> QualType.isPtr() {
    return this.rawType.isPtr();
}

/**
 * Check if the underlying type is a pointer to a certain super type
 *
 * @param superType Super type
 * @return Pointer to super type or not
 */
public f<bool> QualType.isPtrTo(SuperType superType) {
    if !this.isPtr() { return false; }
    const QualType contained = this.getContained();
    return contained.is(superType);
}

/**
 * Check if the underlying type is a reference
 *
 * @return Reference or not
 */
public f<bool> QualType.isRef() {
    return this.rawType.isRef();
}

/**
 * Check if the underlying type is a reference to a certain super type
 *
 * @param superType Super type
 * @return Reference to super type or not
 */
public f<bool> QualType.isRefTo(SuperType superType) {
    if !this.isRef() { return false; }
    const QualType contained = this.getContained();
    return contained.is(superType);
}

/**
 * Check if the underlying type is an array
 *
 * @return Array or not
 */
public f<bool> QualType.isArray() {
    return this.rawType.isArray();
}

/**
 * Check if the underlying type is an array of a certain super type
 *
 * @param superType Super type
 * @return Array of super type or not
 */
public f<bool> QualType.isArrayOf(SuperType superType) {
    if !this.isArray() { return false; }
    const QualType contained = this.getContained();
    return contained.is(superType);
}

/**
 * Check if the underlying type is a const reference
 *
 * @return Const reference or not
 */
public f<bool> QualType.isConstRef() {
    return this.qualifiers.isConst && this.rawType.isRef();
}

/**
 * Check if the current type is an iterator
 *
 * @param node IASTNode
 * @return Iterator or not
 */
public f<bool> QualType.isIterator(const IASTNode* node) {
    // The type must be a struct that implements the iterator interface
    if !this.is(SuperType::TY_STRUCT) { return false; }

    const QualType genericType = QualType(SuperType::TY_GENERIC, String("T"));
    const TypeChainElementData data = TypeChainElementData{/*arraySize=*/ 0u, /*bodyScope=*/ nil<IScope*>, /*hasCaptures=*/ false};
    // ToDo
    return false;
}

/**
 * Check if the current type is an iterable
 * - Arrays are always considered iterable
 * - Otherwise the type must be a struct that implements the iterator interface
 *
 * @param node IASTNode
 * @return Iterable or not
 */
public f<bool> QualType.isIterable(const IASTNode* node) {
    // Arrays are always considered iterable
    if this.isArray() { return true; }
    // Otherwise the type must be a struct that implements the iterator interface
    if !this.is(SuperType::TY_STRUCT) { return false; }

    const QualType genericType = QualType(SuperType::TY_GENERIC, String("T"));
    const TypeChainElementData data = TypeChainElementData{/*arraySize=*/ 0u, /*bodyScope=*/ nil<IScope*>, /*hasCaptures=*/ false};
    //  ToDo
    return false;
}

/**
 * Check if the current type is a string object
 *
 * @return String object or not
 */
public f<bool> QualType.isStringObj() {
    if !this.is(SuperType::TY_STRUCT) { return false; }
    if this.getSubType() != STROBJ_NAME { return false; }
    const IScope* bodyScope = this.getBodyScope();
    const ISourceFile* sourceFile = bodyScope.getSourceFile();
    return sourceFile.isStdFile();
}

/**
 * Check if the current type is an error object
 *
 * @return Error object or not
 */
public f<bool> QualType.isErrorObj() {
    if !this.is(SuperType::TY_STRUCT) { return false; }
    if this.getSubType() != ERROBJ_NAME { return false; }
    const IScope* bodyScope = this.getBodyScope();
    const ISourceFile* sourceFile = bodyScope.getSourceFile();
    return sourceFile.isStdFile();
}

/**
 * Check if the current type has any generic parts
 *
 * @return Generic parts or not
 */
public f<bool> QualType.hasAnyGenericParts() {
    return this.rawType.hasAnyGenericParts();
}

/**
 * Check if copying an instance of the current type would require calling other copy ctors.
 * If this function return true, the type can be copied by calling memcpy.
 *
 * @param node Accessing IASTNode
 * @return Trivially copyable or not
 */
public f<bool> QualType.isTriviallyCopyable(const IASTNode* node) {
    // Heap-allocated values may not be copied via memcpy
    if this.qualifiers.isHeap { return false; }

    // References can't be copied at all
    if this.isRef() { return false; }

    // In case of an array, this item type is determining the copy triviality
    if this.isArray() {
        const QualType baseType = this.getBase();
        return baseType.isTriviallyCopyable();
    }

    // In case of a struct, the member types determine the copy triviality
    if this.is(SuperType::TY_STRUCT) {
        // If the struct has a copy ctor, it is a non-trivially copyable one
        const IStruct* spiceStruct = this.getStruct(node);

        // If the struct itself has a copy ctor, it is not trivially copyable
        const Vector<Arg> args;
        args.pushBack(Arg(this.toConstRef(), false));
        // ToDo
    }

    return true;
}

/**
 * Check if the current type implements the given interface type
 *
 * @param symbolType Interface type
 * @param node Accessing IASTNode
 * @return Struct implements interface or not
 */
public f<bool> QualType.doesImplement(const QualType& implementedInterfaceType, const IASTNode* node) {
    assert this.is(SuperType::TY_STRUCT) && implementedInterfaceType.is(SuperType::TY_INTERFACE);
    const IStruct* spiceStruct = this.getStruct(node);
    assert spiceStruct != nil<IStruct*>;
    // ToDo
    return false;
}

/**
 * Check if a certain input type can be bound (assigned) to the current type->
 *
 * @param inputType Qualified type, which should be bound to the current type
 * @param isTemporary Is the input type a temporary type
 * @return Can be bound or not
 */
public f<bool> QualType.canBind(const QualType& inputType, bool isTemporary) {
    return !isTemporary || inputType.rawType.isRef() || !this.rawType.isRef() || this.isConstRef();
}

/**
 * Check for the matching compatibility of two types.
 * Useful for struct and function matching as well as assignment type validation and function arg matching.
 *
 * @param otherType Type to compare against
 * @param ignoreArraySize Ignore array sizes
 * @param ignoreQualifiers Ignore qualifiers, except for pointer and reference types
 * @param allowConstify Match when the types are the same, but the lhs type is more const restrictive than the rhs type
 * @return Matching or not
 */
public f<bool> QualType.matches(const QualType& otherType, bool ignoreArraySize, bool ignoreQualifiers, bool allowConstify) {
    // Compare type
    if !this.rawType.matches(otherType.rawType, ignoreArraySize) {
        return false;
    }

    // Ignore or compare qualifiers
    return ignoreQualifiers || this.qualifiers.match(otherType.qualifiers, allowConstify);
}

/**
 * Check for the matching compatibility of two types in terms of interface implementation.
 * Useful for function matching as well as assignment type validation and function arg matching.
 *
 * @param structType Type to compare against
 * @return Matching or not
 */
public f<bool> QualType.matchesInterfaceImplementedByStruct(const QualType& structType) {
    if !this.is(SuperType::TY_INTERFACE) || !structType.is(SuperType::TY_STRUCT) {
        return false;
    }

    // Check if the rhs is a struct type that implements the lhs interface type
    const IStruct* spiceStruct = structType.getStruct(nil<ASTNode*>);
    assert spiceStruct != nil<IStruct*>;
    // ToDo
    return true;
}

/**
 * Check if the current type is the same container type as another type.
 * Container types include arrays, pointers, and references.
 *
 * @param other Other type
 * @return Same container type or not
 */
public f<bool> QualType.isSameContainerTypeAs(const QualType& other) {
    return this.rawType.isSameContainerTypeAs(other.rawType);
}

/**
 * Check if the current type is a self-referencing struct type
 *
 * @return Self-referencing struct type or not
 */
public f<bool> QualType.isSelfReferencingStructType(const QualType* typeToCompareWith) {
    if !this.is(SuperType::TY_STRUCT) { return false; }

    // If no type was set by a previous iteration, we set it to the current type
    if typeToCompareWith == nil<const QualType*> {
        typeToCompareWith = this;
    }

    IScope* baseTypeBodyScope = this.getBodyScope();
    for unsigned long i = 0ul; i < baseTypeBodyScope.getFieldCount(); i++ {
        const SymbolTableEntry* field = baseTypeBodyScope.lookupField(i);
        const QualType& fieldType = field.getQualType();
        // Check if the base type of the field matches with the current type, which is also a base type
        // If yes, this is a self-referencing struct type
        if fieldType.getBase() == *typeToCompareWith {
            return true;
        }

        // If the field is a struct, check if it is a self-referencing struct type
        if fieldType.isSelfReferencingStructType(typeToCompareWith) {
            return true;
        }
    }
    return false;
}

/**
 * Check if the given generic type list has a substantiation for the current (generic) type
 *
 * @param genericTypeList Generic type list
 * @return Has substantiation or not
 */
public f<bool> QualType.isCoveredByGenericTypeList(Vector<IGenericType>& genericTypeList) {
    const QualType baseType = this.getBase();
    // Check if the symbol type itself is generic
    if baseType.is(SuperType::TY_GENERIC) {
        // ToDo
    }

    // If the type is non-generic check template types
    bool covered = true;
    // Check template types
    const QualTypeList& baseTemplateTypes = baseType.getTemplateTypes();
    // ToDo

    // If function/procedure, check param and return types
    const dyn options = [SuperType::TY_FUNCTION, SuperType::TY_PROCEDURE];
    if baseType.isOneOf(options, len(options)) {
        const QualTypeList& paramAndReturnTypes = baseType.getFunctionParamAndReturnTypes();
        // ToDo
    }

    return covered;
}

/**
 * Check if the current type needs de-allocation
 *
 * @return Needs de-allocation or not
 */
public f<bool> QualType.needsDeAllocation() {
    if !this.isHeap() { return false; }
    // We only need de-allocation, if we directly point to a heap-allocated type
    // e.g. for heap TestStruct** we don't need to de-allocate, since it is a non-owning pointer to an owning pointer
    return this.isPtr() && !this.isPtrTo(SuperType::TY_PTR);
}

/**
 * Get the name of the symbol type as a string
 *
 * @param name Name stream
 * @param withSize Include the array size for sized types
 * @param ignorePublic Ignore any potential public qualifier
 */
public p QualType.getName(StringStream& name, bool withSize, bool ignorePublic) {
    // Append the qualifiers
    const QualType baseType = this.getBase();
    const TypeQualifiers defaultForSuperType = getTypeQualifiersOf(baseType.getSuperType());
    if !ignorePublic && this.qualifiers.isPublic && !defaultForSuperType.isPublic {
        name << "public ";
    }
    if this.qualifiers.isComposition && !defaultForSuperType.isComposition {
        name << "compose ";
    }
    if this.qualifiers.isConst && !defaultForSuperType.isConst /*ToDo*/ {
        name << "const ";
    }
    if this.qualifiers.isHeap && !defaultForSuperType.isHeap {
        name << "heap ";
    }
    if this.qualifiers.isSigned && !defaultForSuperType.isSigned {
        name << "signed ";
    }
    if this.qualifiers.isUnsigned && !defaultForSuperType.isUnsigned {
        name << "unsigned ";
    }

    // Loop through all chain elements
    this.rawType.getName(name, withSize);
}

/**
 * Get the name of the symbol type as a string
 *
 * @param withSize Include the array size for sized types
 * @param ignorePublic Ignore any potential public qualifier
 * @return Symbol type name
 */
/*public f<String> QualType.getName(bool withSize, bool ignorePublic) {
    StringStream name;
    this.getName(name, withSize, ignorePublic);
    return name.str();
}*/

/**
 * Convert the type to an LLVM type
 *
 * @param sourceFile Source file
 * @return LLVM type
 */
public f<llvm::Type> QualType.toLLVMType(ISourceFile* sourceFile) {
    return this.sourceFile.getLLVMType(this.rawType);
}

/**
 * Retrieve the pointer type to this type
 *
 * @param node ASTNode
 * @return New type
 */
public f<QualType> QualType.toPtr(const ASTNode* node) {
    QualType newType = *this;
    newType.rawType = this.rawType.toPtr(node);
    return newType;
}

/**
 * Retrieve the reference type to this type
 *
 * @param node ASTNode
 * @return New type
 */
public f<QualType> QualType.toRef(const ASTNode* node) {
    QualType newType = *this;
    newType.rawType = this.rawType.toRef(node);
    return newType;
}

/**
 * Retrieve the const reference type of this type
 *
 * @param node ASTNode
 * @return New type
 */
public f<QualType> QualType.toConstRef(const ASTNode* node) {
    QualType newType = this.toRef(node);
    newType.makeConst();
    return newType;
}

/**
 * Retrieve the array type of this type
 *
 * @param node ASTNode
 * @param size Array size
 * @param skipDynCheck Skip dynamic check
 * @return New type
 */
public f<QualType> QualType.toArray(const ASTNode* node, unsigned long size, bool skipDynCheck = false) {
    QualType newType = *this;
    newType.rawType = this.rawType.toArr(newType, size, skipDynCheck);
    return newType;
}

/**
 * Retrieve the non-const type of this type
 *
 * @return New type
 */
public f<QualType> QualType.toNonConst() {
    QualType newType = *this;
    newType.qualifiers.isConst = false;
    return newType;
}

/**
 * Retrieve the contained type of this type
 * This works on pointers, arrays, references and strings (which alias with char*)
 *
 * @return New type
 */
public f<QualType> QualType.getContained() {
    const dyn options = [SuperType::TY_PTR, SuperType::TY_REF, SuperType::TY_ARRAY, SuperType::TY_STRING];
    assert this.isOneOf(options, len(options));
    QualType newType = *this;
    newType.rawType = this.rawType.getContained();
    return newType;
}

/**
 * Retrieve the base type of this type
 *
 * @return New type
 */
public f<QualType> QualType.getBase() {
    QualType newType = *this;
    newType.rawType = this.rawType.getBase();
    return newType;
}

/**
 * Remove reference of this type, if it is a reference
 *
 * @return New type
 */
public f<QualType> QualType.removeReferenceWrapper() {
    return this.isRef() ? this.getContained() : *this;
}

/**
 * Replace the base type with another one
 *
 * @param newBaseType New base type
 * @return The new type
 */
public f<QualType> QualType.replaceBaseType(const QualType& newBaseType) {
    // Create new type
    const IType* newType = this.rawType.replaceBase(newBaseType.getType());
    // Create new qualifiers
    const TypeQualifiers newQualifiers = this.qualifiers.merge(newBaseType.qualifiers);
    // Return the new qualified type
    return QualType(newType, newQualifiers);
}

/**
 * Retrieve the same type, but with lambda captures enabled
 *
 * @return Same type with lambda captures
 */
public f<QualType> QualType.getWithLambdaCaptures(bool enabled = true) {
    // Create new type
    const IType* newType = this.rawType.getWithLambdaCaptures(enabled);
    // Return the new qualified type
    return QualType(newType, this.qualifiers);
}
