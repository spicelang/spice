f<int> main() {
    Lexer lexer = Lexer("./test-file.spice");
    while (!lexer.isEOF()) {
        Token token = lexer.getToken();
        printf("Token: ");
        token.print();
        lexer.advance();
    }
}

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";
import "../../src-bootstrap/ast/ast-nodes";

f<int> main() {
    Lexer lexer = Lexer("./test-file.spice");
    Parser parser = Parser(lexer);
    ASTEntryNode* entryNode = parser.parse();
}*/

/*f<int> main() {
    int i = 123; // Captured by ref
    int j = 321; // Captured by val
    dyn lambda = p() {
        printf("Hello from inside: %d\n", i);
        i++;
        i += j;
        printf("Hello from inside: %d\n", i);
    };
    lambda();
    printf("Hello from outside: %d\n", i);
}*/

/*type Visitable interface {
    p print();
}

type Test1 struct : Visitable {
    int f1
}

p Test1.print() {
    printf("Foo: %d", this.f1);
}

f<int> main() {
    Test1 t1 = Test1{123};
    Visitable* v = &t1;
    v.print();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";

f<int> main() {
    Lexer lexer = Lexer("./file.spice");
    Parser parser = Parser(lexer);
    parser.parse();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "std/time/timer";

f<int> main() {
    Timer timer = Timer();
    timer.start();
    Lexer lexer = Lexer("./file.spice");
    unsigned long i = 1l;
    while (!lexer.isEOF()) {
        Token token = lexer.getToken();
        //printf("Token %d: ", i);
        //token.print();
        lexer.advance();
        i++;
    }
    timer.stop();
    printf("Tokens: %d, Time: %d\n", i, timer.getDurationInMillis());
}*/