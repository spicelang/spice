/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

/*import "std/data/vector" as vector;

f<int> main() {
    dyn v = vector.Vector<int>{};
    v.push(4);
    v.push(2);
}*/

/*import "os-test2" as s1;

f<int> main() {
    s1.Vec v = s1.Vec{11, false};
    v.print();
    //dyn v = s1.Vector<int>{};
    //v.setData<int>(12);
}*/

type TestStruct struct {
    int f1
    int f2
}

f<int> main() {
    TestStruct a = TestStructTypo { 1, 2 };
    printf("Field 1: %d", a.f1);
}