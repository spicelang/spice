import "std/io/filepath";
import "std/os/os";

f<int> main() {
    FilePath path = FilePath("C:\Users\Public\Documents");
    path /= "test.txt";
    assert len(path.toString()) == 34;
    if isWindows() {
        assert path.toString() == "C:\\Users\\Public\\Documents\\test.txt";
    } else {
        assert path.toString() == "C:/Users/Public/Documents/test.txt";
    }
    assert path.getFileName() == "test.txt";
    assert path.getExtension() == "txt";
    assert path.getBaseName() == "test";

    printf("All assertions passed!");
}

/*import "bootstrap/util/block-allocator";
import "bootstrap/util/memory";

f<int> main() {
    DefaultMemoryManager defaultMemoryManager;
    IMemoryManager* memoryManager = &defaultMemoryManager;
    BlockAllocator<int> allocator = BlockAllocator<int>(memoryManager, 10);
}*/