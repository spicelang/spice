import "std/data/unordered-map";
import "std/data/pair";

f<int> main() {
    UnorderedMap<int, String> unorderedMap;

    // Iterate over empty container
    {
        foreach Pair<int&, String&> item : unorderedMap {
            printf("%d: %s\n", item.getFirst(), item.getSecond());
        }
    }

    unorderedMap.upsert(1, String("1"));
    unorderedMap.upsert(2, String("2"));
    unorderedMap.upsert(3, String("3"));
    unorderedMap.upsert(4, String("4"));
    unorderedMap.upsert(5, String("5"));
    unorderedMap.upsert(99, String("99"));
    unorderedMap.upsert(100, String("100"));
    unorderedMap.upsert(1265, String("1265"));
    unorderedMap.upsert(101, String("101"));
    unorderedMap.upsert(102, String("102"));

    // Iterate over filled container
    foreach Pair<int&, String&> item : unorderedMap {
        printf("%d: %s\n", item.getFirst(), item.getSecond());
    }
}


/*f<int> greatestCommonDivisor(int a, int b) {
    while b != 0 {
        int temp = b;
        b = a % b;
        a = temp;
    }
    return a;
}

f<int> main() {
    int a = 56;
    int gcd = greatestCommonDivisor(a, 98);
    printf("GCD of %d and %d is %d.", a, 98, gcd);
}*/