f<int> fibo(int n) {
    printf("Param: %d", n);
    //if n <=1 { return n; }
    //int fibo1 = fibo(n - 1);
    //int fibo2 = fibo(n - 2);
    //return fibo(n - 1) + fibo(n - 2);
    return 0;
}

f<int> main() {
    result = fibo(5);
    printf("%d", result);
    return 0;
}