// Link external functions
ext f<int> pthread_create(byte* /*thread*/, byte* /*attr*/, p() /*start_routine*/, byte* /*arg*/);
ext f<int> pthread_join(byte* /*thread*/, byte** /*retval*/);
ext f<byte*> pthread_self();

public type Thread struct {
    byte* threadId
}

public p Thread.ctor(p() threadRoutine) {
    pthread_create(this.threadId, nil<byte*>, threadRoutine, nil<byte*>);
    //this.threadId = pthread_self();
}

/**
 * Wait synchronous until the thread has terminated
 */
public p Thread.join() {
    pthread_join(this.threadId, nil<byte**>);
}

/**
 * Retrieve the ID of the current thread
 */
public f<byte*> Thread.getId() {
    return this.threadId;
}

/**
 * Retrieve the ID of the current thread
 */
public f<byte*> getThreadId() {
    return pthread_self();
}