import "std/data/pair";

// Generic type definitions
type T dyn;

/**
 * The Iterable interface must be implemented in order to be handled as an iterator by Spice. For instance, all elements,
 * implementing the Iterable interface can be looped over by a standard foreach loop.
 */
public type Iterable<T> interface {
    f<bool> hasNext();
    f<T&> next();
    f<Pair<unsigned long, T&>> nextIdx();
    f<T&> get();
}