f<int> main() {
    thread "non-integer" {
        printf("This is a test");
    }
}