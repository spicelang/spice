import "std/io/cli-parser";

f<int> main(int argc, string[] argv) {
    CliParser cli = CliParser("app-name", "Short description of the app");
    cli.setVersion("v1.0.0");
    cli.setFooter("(c) 2023 by John Doe");

    bool flagValue = false;
    cli.addFlag("--hi", flagValue, "Say Hi");

    cli.parse(argc, argv);

    if flagValue {
        printf("Hi!");
    }
}

/*f<int> main() {
    int z = 2;
    int w = 3;
    p(int&) foo = p(int& x) {
        x += z + w;
    };
    int x = 1;
    foo(x);
    printf("%d", x);
}*/


/*type T int|long;

type TestStruct<T> struct {
    T _f1
    unsigned long length
}

p TestStruct.ctor(const unsigned long initialLength) {
    this.length = initialLength;
}

p TestStruct.printLength() {
    printf("%d\n", this.length);
}

type Alias alias TestStruct<long>;

f<int> main() {
    Alias a = Alias{12345l, (unsigned long) 54321l};
    a.printLength();
    dyn b = Alias(12l);
    b.printLength();
}*/

/*type TestStruct struct {
    long lng
    String str
    int i
}

p TestStruct.dtor() {}

f<TestStruct> fct(int& ref) {
    TestStruct ts = TestStruct{ 6l, String("test string"), ref };
    return ts;
}

f<int> main() {
    int test = 987654;
    const TestStruct res = fct(test);
    printf("Long: %d\n", res.lng);
    printf("String: %s\n", res.str.getRaw());
    printf("Int: %d\n", res.i);
}*/