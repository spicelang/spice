public type DeferredLogic struct {
    p() deferredFunc
    bool triggerOnDestruct
    bool alreadyExecuted = false
}

public p DeferredLogic.ctor(p() deferredFunc, bool triggerOnDestruct = true) {
    this.deferredFunc = deferredFunc;
    this.triggerOnDestruct = triggerOnDestruct;
}

public p DeferredLogic.dtor() {
    if this.triggerOnDestruct && !this.alreadyExecuted {
        p() func = this.deferredFunc;
        func();
    }
}

public p DeferredLogic.execute() {
    p() func = this.deferredFunc;
    func();
    this.alreadyExecuted = true;
}

#[test, test.name="Deferred logic"]
public f<bool> testDeferredLogic() {
    int i = 0;
    int j = 1;
    {
        DeferredLogic _ = DeferredLogic(p() {
            printf("Increment!\n");
            //i++;
            //j++;
            printf("i: %d\n", i);
            printf("j: %d\n", j);
        });
        assert i == 0;
    }
    printf("%d\n", i);
    assert i == 1;

    return true;
}
