import "std/runtime/iterator_rt";

f<int> main() {
    int[7] intArray = { 1, 5, 4, 0, 12, 12345, 9 };
    foreach long index, int item : iterate(intArray, len(intArray)) {
        printf("Item for index %d, %d\n", index, item);
    }
}