public const string GLOBAL = "This is a test";