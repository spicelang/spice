// Imports
import "../reader/code-loc";

// Enums
public type TokenType enum {
    INVALID = 0,
    // Keyword tokens
    TYPE_DOUBLE = 1,
    TYPE_INT = 2,
    TYPE_SHORT = 3,
    TYPE_LONG = 4,
    TYPE_BYTE = 5,
    TYPE_CHAR = 6,
    TYPE_STRING = 7,
    TYPE_BOOL = 8,
    TYPE_DYN = 9,
    CONST = 10,
    SIGNED = 11,
    UNSIGNED = 12,
    INLINE = 13,
    PUBLIC = 14,
    HEAP = 15,
    COMPOSE = 16,
    F = 17,
    P = 18,
    IF = 19,
    ELSE = 20,
    SWITCH = 21,
    CASE = 22,
    DEFAULT = 23,
    ASSERT = 24,
    FOR = 25,
    FOREACH = 26,
    DO = 27,
    WHILE = 28,
    IMPORT = 29,
    BREAK = 30,
    CONTINUE = 31,
    FALLTHROUGH = 32,
    RETURN = 33,
    AS = 34,
    STRUCT = 35,
    INTERFACE = 36,
    TYPE = 37,
    ENUM = 38,
    OPERATOR = 39,
    ALIAS = 40,
    UNSAFE = 41,
    NIL = 42,
    MAIN = 43,
    PRINTF = 44,
    SIZEOF = 45,
    ALIGNOF = 46,
    LEN = 47,
    PANIC = 48,
    EXT = 49,
    TRUE = 50,
    FALSE = 51,
    // Operator tokens
    LBRACE = 52,
    RBRACE = 53,
    LPAREN = 54,
    RPAREN = 55,
    LBRACKET = 56,
    RBRACKET = 57,
    LOGICAL_OR = 58,
    LOGICAL_AND = 59,
    BITWISE_OR = 60,
    BITWISE_XOR = 61,
    BITWISE_AND = 62,
    PLUS_PLUS = 63,
    MINUS_MINUS = 64,
    PLUS_EQUAL = 65,
    MINUS_EQUAL = 66,
    MUL_EQUAL = 67,
    DIV_EQUAL = 68,
    REM_EQUAL = 69,
    SHL_EQUAL = 70,
    SHR_EQUAL = 71,
    AND_EQUAL = 72,
    OR_EQUAL = 73,
    XOR_EQUAL = 74,
    PLUS = 75,
    MINUS = 76,
    MUL = 77,
    DIV = 78,
    REM = 79,
    NOT = 80,
    BITWISE_NOT = 81,
    GREATER = 82,
    LESS = 83,
    GREATER_EQUAL = 84,
    LESS_EQUAL = 85,
    SHL = 86,
    SHR = 87,
    EQUAL = 88,
    NOT_EQUAL = 89,
    ASSIGN = 90,
    QUESTION_MARK = 91,
    SEMICOLON = 92,
    COLON = 93,
    COMMA = 94,
    DOT = 95,
    ARROW = 96,
    SCOPE_ACCESS = 97,
    ELLIPSIS = 98,
    FCT_ATTR_PREAMBLE = 99,
    MOD_ATTR_PREAMBLE = 100,
    // Regex tokens
    DOUBLE_LIT = 101,
    INT_LIT = 102,
    SHORT_LIT = 103,
    LONG_LIT = 104,
    CHAR_LIT = 105,
    STRING_LIT = 106,
    IDENTIFIER = 107,
    TYPE_IDENTIFIER = 108,
    // Skipped tokens
    DOC_COMMENT = 109,
    BLOCK_COMMENT = 110,
    LINE_COMMENT = 111,
    EOF = 112
}

public type Token struct {
    public TokenType tokenType
    public String text
    public CodeLoc codeLoc
}

public p Token.ctor(TokenType tokenType) {
    this.tokenType = tokenType;
}

public p Token.ctor(TokenType tokenType, String text, const CodeLoc& codeLoc) {
    this.tokenType = tokenType;
    this.text = text;
    this.codeLoc = codeLoc;
}

public p Token.ctor(TokenType tokenType, string text, const CodeLoc& codeLoc) {
    this.ctor(tokenType, String(text), codeLoc);
}

public p Token.print() {
    printf("Token(type=%d, text=\"%s\", line=%d, col: %d)\n", this.tokenType, this.text, this.codeLoc.line, this.codeLoc.col);
}