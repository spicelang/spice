import "std/io/cli-parser";
import "std/text/print";

type CliOptions struct {
    bool sayHi = false
}

p callback(bool& value) {
    printf("Callback called with value %d\n", value);
}

f<int> main(int argc, string[] argv) {
    // Setup simple cli
    CliParser cli = CliParser("spice", "This is a test tool");
    cli.setVersion("0.1.0");
    cli.setFooter("(c) Marc Auberer 2023");

    // Setup cli flags
    CliOptions options;
    cli.addFlag("--hi", options.sayHi, "Say hi to the user");
    cli.addFlag("--callback", callback, "Call a callback function");
    cli.addFlag("-cb", p(bool& value) {
        printf("CB called with value %d\n", value);
    }, "Call a callback function");

    // Parse cli arguments
    cli.parse(argc, argv);

    // Print hi if requested
    if options.sayHi {
        println("Hi!");
    }
}

/*f<int> main() {
    int z = 2;
    int w = 3;
    p(int&) foo = p(int& x) {
        x += z + w;
    };
    int x = 1;
    foo(x);
    printf("%d", x);
}*/


/*type T int|long;

type TestStruct<T> struct {
    T _f1
    unsigned long length
}

p TestStruct.ctor(const unsigned long initialLength) {
    this.length = initialLength;
}

p TestStruct.printLength() {
    printf("%d\n", this.length);
}

type Alias alias TestStruct<long>;

f<int> main() {
    Alias a = Alias{12345l, (unsigned long) 54321l};
    a.printLength();
    dyn b = Alias(12l);
    b.printLength();
}*/

/*type TestStruct struct {
    long lng
    String str
    int i
}

p TestStruct.dtor() {}

f<TestStruct> fct(int& ref) {
    TestStruct ts = TestStruct{ 6l, String("test string"), ref };
    return ts;
}

f<int> main() {
    int test = 987654;
    const TestStruct res = fct(test);
    printf("Long: %d\n", res.lng);
    printf("String: %s\n", res.str.getRaw());
    printf("Int: %d\n", res.i);
}*/