import "std/type/type-conversion";

f<int> main() {
    printf("Result: %d\n", toInt(true));
}