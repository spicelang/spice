type T dyn;

type Optional<T> struct {}

p Optional.ctor() {}

f<int> main() {
     dyn oi = Optional();
}