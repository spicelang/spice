f<int> test(string _input) {
    return 12;
}

f<int> invoke(f<int>(string) fctPtr) {
    return fctPtr("string");
}

f<int> main() {
    f<int>(string) testFct = test;
    int i = invoke(testFct);
    printf("%d", i);
}