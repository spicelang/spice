f<int> dummy() {
    return 0;
}