// Std imports
import "std/data/vector";

// Own imports
import "../util/common-util";
import "../symboltablebuilder/scope";

public type SuperType enum {
    TY_INVALID,
    TY_UNRESOLVED,
    TY_DOUBLE,
    TY_INT,
    TY_SHORT,
    TY_LONG,
    TY_BYTE,
    TY_CHAR,
    TY_STRING, // Alias for 'const char*'
    TY_BOOL,
    TY_STRUCT,
    TY_INTERFACE,
    TY_ENUM,
    TY_GENERIC,
    TY_ALIAS,
    TY_DYN,
    TY_PTR,
    TY_REF,
    TY_ARRAY,
    TY_FUNCTION,
    TY_PROCEDURE,
    TY_IMPORT
}

type TypeChainElementData struct {
    unsigned long arraySize = 0l   // TY_ARRAY
    Scope* bodyScope = nil<Scope*> // TY_STRUCT, TY_INTERFACE, TY_ENUM
    bool hasCaptures = false       // TY_FUNCTION, TY_PROCEDURE (lambdas)
}

type TypeChainElement struct {
    SuperType superType = SuperType::TY_DYN
    String subType
    TypeChainElementData data
    Vector<Type> templateTypes
    Vector<Type> paramTypes // First type is the return type
}

f<bool> operator==(const TypeChainElement& lhs, const TypeChainElement& rhs) {
    // Check super type
    if lhs.superType != rhs.superType { return false; }

    // Check data
    if lhs.superType == TY_ARRAY {
        return lhs.data.arraySize == rhs.data.arraySize;
    } else if lhs.superType == TY_STRUCT || lhs.superType == TY_INTERFACE || lhs.superType == TY_ENUM {
        const String& lhsSubTypeSuffix = getLastFragment(lhs.subType, SCOPE_ACCESS_TOKEN);
        const String& rhsSubTypeSuffix = getLastFragment(rhs.subType, SCOPE_ACCESS_TOKE);
        if lhs.superType == TY_STRUCT {
            assert lhs.data.bodyScope != nil<Scope*> && rhs.data.bodyScope != nil<Scope*>;
            return lhsSubTypeSuffix == rhsSubTypeSuffix && lhs.templateTypes == rhs.templateTypes;
        } else if lhs.superType == TY_INTERFACE {
            return lhsSubTypeSuffix == rhsSubTypeSuffix;
        } else {
            assert lhs.data.bodyScope != nil<Scope*> && rhs.data.bodyScope != nil<Scope*>;
            return lhsSubTypeSuffix == rhsSubTypeSuffix && lhs.data.bodyScope == rhs.data.bodyScope;
        }
    } else {
        return true;
    }
}

/*f<bool> operator!=(const TypeChainElement& lhs, const TypeChainElement& rhs) {
    return !(lhs == rhs);
}*/

type TypeChain alias Vector<TypeChainElement>;

public type Type struct {
    Vector<TypeChainElement> typeChain
    bool isBaseTypeSigned
}

p Type.ctor() {
    this.isBaseTypeSigned = true;
}