public type IType interface {

}