type UnusedStruct struct {}

f<int> main() {}