type Person struct {
    string firstName
    string lastName
    unsigned int age
}

p birthday(Person* person) {
    person.age++;
}

f<int> main() {
    dyn mike = Person { "Mike", "Miller", 32u };
    printf("Person: %s, %s\n", mike.lastName, mike.firstName);
    printf("Age before birthday: %d\n", mike.age);
    birthday(&mike);
    printf("Age after birthday: %d\n", mike.age);
}