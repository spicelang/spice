import "std/data/vector";
import "std/data/linked-list";
import "std/runtime/iterator_rt";
import "std/data/pair";
import "std/math/hash";

// Generic types for key and value
type K dyn;
type V dyn;

public type HashTable<K, V> struct {
    Vector<LinkedList<Pair<K, V>>> table
    unsigned long bucketCount
}

public p HashTable.ctor(unsigned long bucketCount = 1000l) {
    this.bucketCount = bucketCount;
}

public p HashTable.insert(const K& key, const V& value) {
    const unsigned long index = hash(key);
    foreach dyn bucket : iterate(this.table) {
        if bucket.getFirst() == key {
            bucket.add(Pair<K, V>(key, value));
            return;
        }
    }
    this.table.pushBack(LinkedList<Pair<K, V>>());
    LinkedList<Pair<K, V>>& bucket = this.table.back();
    bucket.add(Pair<K, V>(key, value));
}

public p HashTable.delete(const K& key) {
    const unsigned long index = hash(key);
    const LinkedList<Pair<K, V>>& bucket = this.table.at(index);

    for unsigned long i = 0l; i < bucket.getSize(); i++ {
        Pair<K, V>& candidate = bucket.at(i);
        if candidate.getFirst() == key {
            bucket.remove(i);
            return;
        }
    }
}

public f<V*> HashTable.search(const K& key) {
    unsigned long index = hash(key);
    const LinkedList<Pair<K, V>>& bucket = this.table.at(index);

    for unsigned long i = 0l; i < bucket.getSize(); i++ {
        Pair<K, V>& candidate = bucket.at(i);
        if candidate.getFirst() == key {
            return &candidate.getSecond();
        }
    }
    return nil<V*>;
}