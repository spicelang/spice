f<string> getOsName() {
    return "linux";
}