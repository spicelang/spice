type T dyn;

type Vec struct {
    T genericField
}

f<int> main() {
    Vec v = Vec{};
}