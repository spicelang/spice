// TEST: --sanitizer=thread -g

import "std/os/thread";

int COUNTER = 0;

p worker() {
    for int i = 0; i < 1000000; i++ {
        COUNTER++;
    }
}

f<int> main() {
    Thread thread1 = Thread(worker);
    Thread thread2 = Thread(worker);
    thread1.run();
    thread2.run();
    thread1.join();
    thread2.join();
}