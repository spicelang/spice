import "source2";

public type Car struct : Driveable {
    bool driving
}

p Car.ctor() {
    this.driving = false;
}

p Car.drive(int _param) {
    this.driving = true;
}

f<bool> Car.isDriving() {
    return this.driving;
}

f<int> main() {
    Car car = Car();
    Driveable* driveable = &car;
    driveable.drive(12);
    printf("Is driving: %d", driveable.isDriving());
}