public const int ANONYMOUS = -1;