f<int> main() {
    int val = 1;
    val += ((1++)--) * 2 << 2;
    printf("Value: %d\n", val);
}