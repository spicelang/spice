import "std/io/csv";

f<int> main() {
    CSVParser parser = CSVParser("test.csv");

}