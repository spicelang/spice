type NotAPointer struct {}

f<int> main() {
    NotAPointer nonPtr = NotAPointer {};
    printf("%p", nonPtr);
}