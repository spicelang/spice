import "std/time/timer";
import "std/time/delay";

f<bool> isInRange(unsigned long duration, unsigned long expectedDuration, unsigned int delta) {
    printf("Check for %d +/-%d, got %d\n", expectedDuration, delta, duration);
    return duration >= expectedDuration - delta && duration <= expectedDuration + delta;
}

f<int> main() {
    // Normal start/stop scenario
    Timer t = Timer();
    assert t.getDuration() == 0l;
    t.start();
    delay(10);
    t.stop();
    assert isInRange(t.getDuration(), 10l, 3); // 10 +/-3 millis

    // Start/pause/resume/stop with seconds
    unsigned long duration = 0l;
    t = Timer(TimerMode::MICROS, &duration);
    assert t.getDuration() == 0l;
    assert duration == 0l;
    t.start();
    delay(10);
    t.pause();
    delay(100);
    t.resume();
    delay(10);
    t.stop();
    assert isInRange(duration, 20000l, 5000); // 20000 +/-5000 micros

    printf("All assertions passed");
}