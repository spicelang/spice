import "std/io/cli-option";
import "std/runtime/iterator_rt";
import "std/os/os";

// Generic types
type T bool|string|int|long|short;

public type CliParser struct {
    string appName
    string appDescription
    string footer
    string versionString
    //Vector<CliOption> options
    Vector<CliOption<bool>> flags
    bool allowUnknownOptions = false
}

public p CliParser.ctor(string appName, string appDescription = "") {
    this.appName = appName;
    this.appDescription = appDescription;
    //this.options = Vector<CliOption>();
    this.flags = Vector<CliOption<bool>>();
}

public p CliParser.setVersion(string versionString) {
    this.versionString = versionString;
}

public p CliParser.setFooter(string footer) {
    this.footer = footer;
}

public p CliParser.allowUnknownOptions() {
    this.allowUnknownOptions = true;
}

public p CliParser.addOption<T>(string name, T& targetVariable, string description) {
    //const CliOption option = CliOption<T>(name, targetVariable, description);
    //this.options.pushBack(option);
}

public p CliParser.addFlag(string name, bool& targetVariable, string description) {
    const dyn flag = CliOption<bool>(name, targetVariable, description);
    this.flags.pushBack(flag);
}

public p CliParser.addFlag(string name, p(bool&) callback, string description) {
    const dyn flag = CliOption<bool>(name, callback, description);
    this.flags.pushBack(flag);
}

public f<int> CliParser.parse(unsigned int argc, string[] argv) {
    for unsigned int argNo = 1; argNo < argc; argNo++ {
        const string arg = argv[argNo];

        // Check all commonly used flags
        if (arg == "-v" || arg == "--version") { // Version info
            this.printVersion();
            return EXIT_CODE_SUCCESS;
        }
        if (arg == "-h" || arg == "--help") { // Help
            this.printHelp(argv[0]);
            return EXIT_CODE_SUCCESS;
        }

        // Check for flags
        foreach const CliOption<bool>& flag : iterate(this.flags) {
            if (arg == flag.getName()) {
                flag.setToTrue();
                flag.callCallback(true);
                continue 2; // Continue with next argument
            }
        }

        // We could not match the argument
        if !this.allowUnknownOptions {
            printf("Unknown argument: %s\n", arg);
            return EXIT_CODE_ERROR;
        }
    }
    return EXIT_CODE_SUCCESS; // Parsing was successful, return success exit code
}

p CliParser.printHelp(string fileName) {
    printf("%s\n\nUsage: %s [options]\n\nFlags:\n", this.appDescription, fileName);
    foreach const CliOption<bool>& flag : iterate(this.flags) {
        printf("%s\t\t\t%s\n", flag.getName(), flag.getDescription());
    }
    printf("\n%s\n", this.footer);
}

p CliParser.printVersion() {
    printf("%s\n", this.versionString);
}