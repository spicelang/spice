needs_ext malloc(int);
needs_ext free(char*);
needs_ext memcpy(char*, char* int);

type String struct {
    char[] value
    int len
    int maxLen
    int growthFactor
}

p String.constructor() {
    this.value = null;
    this.len = 0;
    this.maxLen = 0;
    this.growthFactor = 2;
}

p String.destructor() {
    if this.value != null {
        // Free the allocated heap space
        free(this.value);
    }
}

p String.resize(int newLen) {
    char* newAddr = malloc(newLen);
    char* oldAddr = this.value;
    int len = this.length;
    memcpy(newAddr, oldAddr, len);
    free(oldAddr);
    this.value = newAddr;
    this.maxLen = newLen;
}

p String.appendChar(char c) {
    int len = this.length;
    int maxLen = this.maxLen;

    if len == maxLen { // Sting needs to be grown
        int newMaxLen = maxLen * this.growthFactor;
        this.resize(newMaxLen);
    }

    this.value[length] = c;
    this.len++;
}

p String.clear() {
    this.value = null;
    this.len = 0;
    this.maxLen = 0;
}

f<string> concat(string a, string b) {
    // Return b if a is empty
    int aLen = len(a);
    if aLen == 0 { return b; }

    // Return a if b is empty
    int bLen = len(b);
    if bLen == 0 { return a; }
    
    // Create a new string
    int size = aLen + bLen;
    result = "";
    foreach int pos, char n : a {
        result[pos] = n;
    }
    foreach int pos, char n : b {
        result[aLen + pos] = n;
    }

    return result;
}