import "std/type/byte";

f<int> main() {
    // toDouble()
    double asDouble = toDouble(cast<byte>(15));
    assert asDouble == 15.0;

    // toInt()
    int asInt = toInt(cast<byte>(9));
    assert asInt == 9;

    // toShort()
    short asShort = toShort(cast<byte>(6));
    assert asShort == 6s;

    // toLong()
    long asLong = toLong(cast<byte>(63));
    assert asLong == 63l;

    // toString()
    String asString = toString(cast<byte>(13));
    assert asString.getRaw() == "13";

    // toBool()
    bool asBool1 = toBool(cast<byte>(1));
    assert asBool1 == true;
    bool asBool2 = toBool(cast<byte>(0));
    assert asBool2 == false;

    printf("All assertions succeeded");
}