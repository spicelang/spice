f<int> main() {
    string test = "Hello World!";
    string* testPtr = &test;
    printf("Value1: %s, pointer: %p, value: %s", test, testPtr, *testPtr);
}