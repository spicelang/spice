// Std imports
import "std/data/vector";
import "std/io/filepath";

// Own imports
import "bootstrap/driver";

public type ExternalLinkerInterface struct {
    CliOptions& cliOptions
    Vector<FilePath> objectFilePaths
    Vector<String> linkerFlags
    FilePath outputPath
    bool linkLibMath = false
}

public p ExternalLinkerInterface.ctor(CliOptions& cliOptions) {
    this.cliOptions = cliOptions;
    this.outputPath = cliOptions.outputPath;
}

public p ExternalLinkerInterface.prepare() {
    // Set target to linker
    this.addLinkerFlag("--target=" + this.cliOptions.targetTriple);

    // Static linking
    if this.cliOptions.staticLinking {
        this.addLinkerFlag("-static");
    }

    // Stripping symbols
    if !this.cliOptions.generateDebugInfo {
        this.addLinkerFlag("-Wl,-s");
    }

    switch this.cliOptions.instrumentation.sanitizer {
        case Sanitizer::ADDRESS: {
            this.addLinkerFlag("-lasan");
        }
        case Sanitizer::THREAD: {
            this.addLinkerFlag("-ltsan");
        }
        case Sanitizer::MEMORY: {
            this.addLinkerFlag("-L$(clang -print-resource-dir)/lib/x86_64-unknown-linux-gnu");
            this.addLinkerFlag("-lclang_rt.msan");
            this.requestLibMathLinkage();
        }
        case Sanitizer::TYPE: {
            this.addLinkerFlag("-L$(clang -print-resource-dir)/lib/x86_64-unknown-linux-gnu");
            this.addLinkerFlag("-lclang_rt.tysan");
        }
    }

    // Web Assembly
    if this.cliOptions.targetArch == TARGET_WASM32 || this.cliOptions.targetArch == TARGET_WASM64 {
        this.addLinkerFlag("-nostdlib");
        this.addLinkerFlag("-Wl,--no-entry");
        this.addLinkerFlag("-Wl,--export-all");
    }
}

/**
 * Start the linking process
 */
public p ExternalLinkerInterface.link() {

    // ToDo
}

/**
 * Add another object file to be linked when calling 'link()'
 *
 * @param objectFilePath Path to the object file
 */
public p ExternalLinkerInterface.addObjectFilePath(const FilePath& objectFilePath) {
    this.objectFilePaths.pushBack(objectFilePath);
}

/**
 * Add another linker flag for the call to the linker executable
 *
 * @param linkerFlag Linker flag
 */
public p ExternalLinkerInterface.addLinkerFlag(string linkerFlag) {
    this.linkerFlags.pushBack(String(linkerFlag));
}

/**
 * Add another linker flag for the call to the linker executable
 *
 * @param linkerFlag Linker flag
 */
public p ExternalLinkerInterface.addLinkerFlag(const String& linkerFlag) {
    this.linkerFlags.pushBack(linkerFlag);
}

/**
 * Add another source file to compile and link in (C or C++)
 *
 * @param additionalSource Additional source file
 */
public p ExternalLinkerInterface.addAdditionalSourcePath(FilePath additionalSource) {
    // Check if the file exists
    if !additionalSource.exists() {
        const String msg = "The additional source file '" + additionalSource.toGenericString() + "' does not exist";
        panic(Error(msg.getRaw()));
    }

    // Add the file to the linker
    this.addObjectFilePath(additionalSource);
}

/**
 * Link against libmath a.k.a. -lm
 */
public p ExternalLinkerInterface.requestLibMathLinkage() {
    this.linkLibMath = true;
}
