// Std imports
import "std/type/Any" as any;
import "std/data/Vector" as vec;
import "std/type/long" as longTy;

// Own imports
import "AbstractAstVisitor" as vis;
import "../util/CodeLoc" as codeclLoc;
import "../symbol/SymbolType" as st;

/**
 * Saves a constant value for an AST node to realize features like array-out-of-bounds checks
 */
public type CompileTimeValue struct {
    double doubleValue
    int intValue
    short shortValue
    long longValue
    byte byteValue
    char charValue
    char *stringValue
    bool boolValue
}

public type Visitable interface {
    f<any::Any> accept(vis::AbstractAstVisitor*);
}

// =========================================================== AstNode ===========================================================

public type AstNode struct : Visitable {
    AstNode* parent
    vec::Vector<AstNode*> children
    const cl::CodeLoc codeLoc
    string errorMessage
    unsigned long manIdx
    vec::Vector<symbolType::SymbolType> symbolTypes
    CompileTimeValue compileTimeValue
    string compileTimeStringValue
    bool hasDirectCompileTimeValue
}

p AstNode.ctor(AstNode *parent, cl::CodeLoc codeLoc) {
    this.parent = parent;
    this.codeLoc = codeLoc;
    this.manIdx = longTy::MAX_VALUE;
    this.hasDirectCompileTimeValue = false;
}

public f<any::Any> AstNode.accept(vis::AbstractAstVisitor* _) {
    assert false; // Please override at child level
}

// ========================================================== EntryNode ==========================================================

public type AstEntryNode struct : Visitable {
    AstNode astNode
}

public p AstEntryNode.ctor() {

}