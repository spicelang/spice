f<int> main() {
    String strA = String("Hello ");
    String strB = String("World!");
    //String strC = strA + strB;
    printf("%d", strA);
    printf("%d", strB);
    //printf("%d", strC);
}