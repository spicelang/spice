import "std/text/analysis";

// Constants
const int ASCII_SHIFT_OFFSET = 32;
const int MIN_LOWER_CHAR = 97;
const int MAX_LOWER_CHAR = 122;
const int MIN_UPPER_CHAR = 65;
const int MAX_UPPER_CHAR = 90;

/**
 * Returns a formatted storage string (e.g. 1.4 MB for 1,500,000)
 *
 * @return Formatted size string
 */
public f<String> formatStorageSize(long bytes) {
    // ToDo when string concatenation works
    return String("");
}

/**
 * Returns the given text in caps
 *
 * @return Text in caps
 */
/*public p toUpper(String& text) {
    foreach char& c : text {
        if c >= (char) MIN_LOWER_CHAR && c <= (char) MAX_LOWER_CHAR {
            c += (char) ASCII_SHIFT_OFFSET;
        }
    }
    return text;
}*/

/**
 * Returns the given char as upper case version
 *
 * @return Char in upper case
 */
public f<char> toUpper(char c) {
    if c >= (char) MIN_LOWER_CHAR && c <= (char) MAX_LOWER_CHAR {
        c += (char) ASCII_SHIFT_OFFSET;
    }
    return c;
}

/**
 * Returns the given text in all-lower letters
 *
 * @return Text in all-lower letters
 */
/*public p toLower(String& text) {
    foreach char& c : text {
        if c >= (char) MIN_UPPER_CHAR && c <= (char) MAX_UPPER_CHAR {
            c -= ASCII_SHIFT_OFFSET;
        }
    }
    return text;
}*/

/**
 * Returns the given char as lower case version
 *
 * @return Char in lower case
 */
public f<char> toLower(char c) {
    if c >= (char) MIN_UPPER_CHAR && c <= (char) MAX_UPPER_CHAR {
        c -= (char) ASCII_SHIFT_OFFSET;
    }
    return c;
}

/**
 * Returns the given text in capitalized form
 *
 * @return Capitalized text
 */
/*public p capitalize(String& text) {
    if text[0] >= (char) MIN_LOWER_CHAR && text[0] <= (char) MAX_LOWER_CHAR {
        text[0] += (char) ASCII_SHIFT_OFFSET;
    }
    return text;
}*/

/**
 * Returns the trimmed string of the given text
 *
 * @return Trimmed string
 */
/*public f<String> trim(const String& input) {
    unsigned long start = 0l;
    unsigned long end = input.getLength() - 1l;

    while isWhitespace(input[start]) {
        start++;
    }
    while isWhitespace(input[end]) {
        end--;
    }

    return input.substring(start, end);
}*/