// Constants
const unsigned long INITIAL_ALLOC_COUNT = 5l;
const unsigned int RESIZE_FACTOR = 2;

// Link external functions
ext<byte*> malloc(long);
ext<byte*> realloc(byte*, int);
ext free(byte*);
ext<byte*> memcpy(byte*, byte*, int);

// Add generic type definition
type T dyn;

/**
 * A vector in Spice is a commonly used data structure, which can be used to represent a list of items.
 *
 * Time complexity:
 * Insert: O(1)
 * Delete: O(n * m); n = deleted elements, m = moved elements
 * Search: O(n)
 *
 * Vectors pre-allocate space using an initial size and a resize factor to not have to re-allocate
 * with every item pushed.
 */
public type Vector<T> struct {
    T* contents             // Pointer to the first data element
    unsigned long capacity  // Allocated number of items
    unsigned long size      // Current number of items
    unsigned int itemSize   // Size of a single item
}

public p Vector.ctor(unsigned int initAllocItems) {
    this.ctor((long) initAllocItems);
}

public p Vector.ctor(unsigned long initAllocItems = INITIAL_ALLOC_COUNT) {
    // Allocate space for the initial number of elements
    this.itemSize = sizeof(type T) / 8;
    unsafe {
        this.contents = (T*) malloc(this.itemSize * initAllocItems);
    }
    this.size = 0l;
    this.capacity = initAllocItems;
}

public p Vector.ctor(unsigned long initAllocItems, const T& defaultValue) {
    // Allocate space for the initial number of elements
    this.ctor(initAllocItems);
    // Fill in the default values
    for int index = 0; index < initAllocItems; index++ {
        unsafe {
            this.contents[index] = defaultValue;
        }
    }
    this.size = initAllocItems;
}

public p Vector.dtor() {
    // Free all the memory
    unsafe {
        free((byte*) this.contents);
    }
}

/**
 * Checks if the vector contains any items at the moment
 *
 * @return Empty or not empty
 */
public f<bool> Vector.isEmpty() {
    return this.size == 0;
}

/**
 * Checks if the vector exhausts its capacity and needs to resize at the next call of push
 *
 * @return Full or not full
 */
public f<bool> Vector.isFull() {
    return this.size == this.capacity;
}

/**
 * Add an item at the end of the vector
 */
public p Vector.pushBack<T>(const T& item) {
    // Check if we need to re-allocate memory
    if this.isFull() {
        this.resize(this.capacity * RESIZE_FACTOR);
    }

    // Insert the element at the back
    unsafe {
        this.contents[(int) this.size++] = item;
    }
}

/**
 * Get an item at a certain index
 *
 * @return item at index
 */
public f<T&> Vector.get(unsigned long index) {
    assert index < this.size;
    unsafe {
        return this.contents[index];
    }
}

/**
 * Get an item at a certain index
 *
 * @return item at index
 */
public f<T&> Vector.get(unsigned int index) {
    return this.get((unsigned long) index);
}

/**
 * Removes all items from the vector
 */
public p Vector.clear() {
    this.size = 0l;
}

/**
 * Reserves `itemCount` items
 */
public p Vector.reserve(unsigned long itemCount) {
    if itemCount > this.capacity {
        this.resize(itemCount);
    }
}

/**
 * Reserves `itemCount` items
 */
public p Vector.reserve(unsigned int itemCount) {
    if itemCount > this.capacity {
        this.resize((long) itemCount);
    }
}

/**
 * Retrieve the current size of the vector
 *
 * @return Current size of the vector
 */
public f<long> Vector.getSize() {
    return this.size;
}

/**
 * Retrieve the current capacity of the vector
 *
 * @return Current capacity of the vector
 */
 public f<long> Vector.getCapacity() {
     return this.capacity;
 }

/**
 * Frees allocated memory that is not used by the queue
 */
public p Vector.pack() {
    // Return if no packing is required
    if this.isFull() { return; }
    // Pack the array
    this.resize(this.size);
}

/**
 * Re-allocates heap space for the queue contents
 */
p Vector.resize(unsigned long itemCount) {
    // Allocate the new memory
    unsafe {
        byte* oldAddress = (byte*) this.contents;
        int newSize = (int) (this.itemSize * itemCount);
        T* newMemory = (T*) realloc(oldAddress, newSize);
        this.contents = newMemory;
    }
    // Set new capacity
    this.capacity = itemCount;
}