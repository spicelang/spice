//import "std/type/int" as unused;

import "os-test2" as s1;

f<int> main() {
    dyn v = s1::Vector<int>{};
    v.setData(12);
    printf("Data: %d\n", v.data);
    v.setData(1.5);
    printf("Data: %d\n", v.data);
}