f<string> testFunction() {
    return "Hello World!";
}