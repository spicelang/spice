type Letter struct {
    string content
}

f<string> Letter.getContent() {
    return this.content;
}

p Letter.setContent(string text) {
    this.content = text;
}

f<int> main() {
    dyn letter = Letter { "No content" };
    letter.setContent("Hello World!");
    printf("Content: %s\n", letter.getContent());
}

/*import "std/time/timer";
import "../../src-bootstrap/lexer/lexer";

f<int> main(int argc, string[] argv) {
    Timer timer = Timer();
    timer.start();
    Lexer lexer = Lexer(argv[1]);
    unsigned long i = 1l;
    while (!lexer.isEOF()) {
        Token token = lexer.getToken();
        //printf("Token %d: ", i);
        //token.print();
        lexer.advance();
        i++;
    }
    timer.stop();
    printf("Tokens: %d in %d ms\n", i, timer.getDurationInMillis());
}*/

/*type Visitable interface {
    p print();
}

type Test1 struct : Visitable {
    int f1
}

p Test1.print() {
    printf("Foo: %d", this.f1);
}

f<int> main() {
    Test1 t1 = Test1{123};
    Visitable* v = &t1;
    v.print();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "../../src-bootstrap/parser/parser";

f<int> main() {
    Lexer lexer = Lexer("./file.spice");
    Parser parser = Parser(lexer);
    parser.parse();
}*/

/*import "../../src-bootstrap/lexer/lexer";
import "std/time/timer";

f<int> main() {
    Timer timer = Timer();
    timer.start();
    Lexer lexer = Lexer("./file.spice");
    unsigned long i = 1l;
    while (!lexer.isEOF()) {
        Token token = lexer.getToken();
        //printf("Token %d: ", i);
        //token.print();
        lexer.advance();
        i++;
    }
    timer.stop();
    printf("Tokens: %d, Time: %d\n", i, timer.getDurationInMillis());
}*/