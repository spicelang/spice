f<int> spawnInteger() {
    return 7;
}