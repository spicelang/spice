type Nested struct {
    string nested1
    bool* nested2
}

type TestStruct struct {
    int* field1
    double field2
    Nested* nested
}

f<int> main() {
    int input = 12;
    bool boolean = true;
    Nested nestedInstance = new Nested { "Hello World!", &boolean };
    dyn instance = new TestStruct { &input, 46.34, &nestedInstance };
    TestStruct instance1 = instance;
    instance1.field2 = 1.123;
}