ext f<dyn> exteralFunction();

f<int> main() {
    extFunction(1, 3);
}