import "std/os/os" as os;

f<int> main() {
    if isLinux() {
        assert os::OS_NAME == "linux";
    } else if isWindows() {
        assert os::OS_NAME == "windows";
    }
}