return 6.7;

f<int> main() {
    printf("Hello world!");
}