#[non.existing.attr = 321]
f<int> main() {
    printf("Do nothing ...");
}