/**
 * A NumberIterator in Spice can be used to iterate over
 */
public type NumberIterator<U> struct : Iterable<U> {
    U lowerBound
    U upperBound
    unsigned long index
}

public p NumberIterator.ctor(U lowerBound, U upperBound) {
    this.lowerBound = lowerBound;
    this.upperBound = upperBound;
    this.index = 0;
}

public inline const f<bool> NumberIterator.hasNext() {
    return this.lowerBound + this.index <= this.upperBound;
}

public inline f<U*> NumberIterator.next() {
    assert this.hasNext();
    this.index++;
    return this.data;
}

public inline f<U&> NumberIterator.get() {
    return this.lowerBound + this.index;
}