// Imports
import "std/type/long";

public type CodeLoc struct {
    unsigned long line
    unsigned long col
    string sourceFilePath
}

public p CodeLoc.ctor(unsigned long line, unsigned long col, string sourceFilePath = "") {
    this.line = line;
    this.col = col;
    this.sourceFilePath = sourceFilePath;
}

/**
 * Returns the code location as a string for using it as a map key or similar
 *
 * @return Code location string
 */
public f<string> CodeLoc.toString() {
    return "L" + toString(this.line) + "C" + toString(this.col);
}

/**
 * Returns the code location in a pretty form
 *
 * @return Pretty code location
 */
public f<String> CodeLoc.toPrettyString() {
    String codeLocStr = String(intTy.toString(line));
    if this.sourceFilePath.empty() {
        return toString(line) + ":" + toString(this.col);
    }
    return this.sourceFilePath + ":" + toString(this.line) + ":" + toString(this.col);
}

/**
 * Returns the line number in a pretty form
 *
 * @return Pretty line number
 */
public f<string> CodeLoc.toPrettyLine() {
    return "l" + toString(this.line);
}
