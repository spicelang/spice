//import "std/iterators/ranges";
import "std/data/vector";
import "std/data/pair";

f<int> main() {
    Vector<Pair<int, string>> pairVector = Vector<Pair<int, string>>();
    pairVector.pushBack(Pair<int, string>(0, "Hello"));
    pairVector.pushBack(Pair<int, string>(1, "World"));

    Pair<int, string> p1 = pairVector.get(1);
    printf("Hello %s!\n", p1.getSecond());

    //NumberIterator<int> it = range(1, 5);
    /*for (
        dyn it = range(1l, 10l);
        it.hasNext();
        it.next()
    ) {
        printf("%d\n", it.get());
    }*/

    /*foreach int i : range(1, 3) {
        printf("%d\n", i);
    }*/
}