/*type StringStruct struct {
    int len
    char* value
    int maxLen
    int growthFactor
}

p StringStruct.appendChar(char c) {
    this.value[1] = c;
}

f<int> main() {
    StringStruct a = StringStruct {};
    a.appendChar('A');
}*/

/*import "std/runtime/string_rt" as str;

f<int> main() {
    str.StringStruct a = str.StringStruct {};
    a.constructor();
    printf("String: %s\n", a.value);
    a.appendChar('A');
    printf("String: %s\n", a.value);
    a.destructor();
}*/

type Person struct {
    string firstName
    string lastName
    int age
}

p birthday(Person* person) {
    person.age++;
}

f<int> main() {
    dyn mike = Person { "Mike", "Miller", 32 };
    printf("Person: %s, %s", mike.lastName, mike.firstName);
    printf("Age before birthday: %d", mike.age);
    birthday(&mike);
    printf("Age after birthday: %d", mike.age);
}